// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HD4TCI+# K./<<'78;J&7_;F0!K@@U M7B=:IOF]%5RY+7S/X3K6#Q@  
HF[8?%I?C;.TMEXKO4>GZ2]F>_#XU05)4<('9!P(AI$:V=8(DV'^6P0  
HL,C3OZTJV"Y*W(#0"7*>3/30^)) EQ^49@L2NL*,$J!ZUMSD39[)%P  
HOZ)4(EP[_!>WT SW<CG1^?"F8?[7Z":\^+'R=_L.F@C)>-9UJ8I4S@  
H &5![T:S1Z=,H)F1B^'0OQ$3KT4CS\SY,&DM<BTCG2H7]>N9&FJ!90  
`pragma protect encoding=(enctype="uuencode",bytes=3728        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@J'X"S <*ZO7(,UA_1*T4=":2MMW1! GWX*41$GY.KA@ 
@^=9'=.*DS3T"*#:[Z>_]AY#>.(2(8W=3Q"JDE*^/H:< 
@^S$&U&@ZDZD>$6C]1J ,T'2"9(ATV:'NL[F?+FPX"&L 
@1;>_Y:(*8"@S?"LJ@63]$*4^^]>IH9^<38?%/TF.]/0 
@KZO*,-Y2JQJGLTF?=V&DH#292$GM9C:3SS,Z/2Q6O=0 
@+?RS+I.76LB,.HNB-XE_W'<:_LK*LA*6[M(BLYM3SRX 
@[UURISSA6#T;I%WL V^4Y"#,V/TR:.K+YS5O(55*A P 
@J#+8:=_7'DQ3@A&7ZF,5?)];LOQ:[$)ZP&U;>Y%60O, 
@UL47(2+0U*#\32)WU&!)*=+F:WD*;_K:+7L2QZT,"HD 
@LV3V@ILW1@AKE(EC V++1-_.%F-;AJMVK=-Z#V9JF?@ 
@@EY<'J"M>"#J,5:< IZOWQ(.[[KN/H0-7K5=#*IS2$8 
@W#!^VR&Q*CG<P-N*CS78RYE) ET<F,-!RM)Q-3 /O-, 
@/_!:8NYC(P/!='T>&VKW2TO!'#RV'_P];V%R"0E'>KX 
@,/ZJ&5U_*T@, &5%58WS)F$'O"N?#+[T5/0Y;\<]XGD 
@-[R2LO/HS>L5([FP4BR*3 &NRYVN;TQ.8"XD7'YU2J  
@Y*5_09P$3Y=X1'@7*,6Q3OFYUV)[/C?KR]T O6).#G0 
@+/L%2<X0M*'M-&R:3U7D)*M@03'+*=6=%B22K1CI *< 
@7#3]4S\=P X_%Q9[5=VVQ($7^_D"WY]B?)IKDBQ543P 
@#F1"+OD9J50!3(Q*I>1<P&?6MMBY&5\SC=@*4 G9Y8T 
@8#TGYC0;:L5;0,4@6&GI=3NX?(T2?8NM>T(FAHE1)AT 
@]7P[LR1L $P>."DTL(5^%;LG+J*EP.?43J0A;(NI]Y\ 
@^QXQ.!U%7-/3'/?6@PE>3Z&IB]4C7\A(:-;S867 @B0 
@_-(\)*UN%NY6*;PW'--M:T])W]@>O@"?S-^:ZM*RQ>4 
@K-?'1M8<\67L>: :[O^T4/YN'I>8[=\91DLC9U;W:'0 
@JEH-M>70*E<H>OYFI.(J,]F3_<^&S:_+)]((1$Z=2OD 
@*1Q[C.VQ*G?:^XIP&6O?3-3D 1*<U!@DI#(BU8GV,8< 
@X=&H]AUBZ0 WGCP!D_@9^XO4RR,]P.Q2MD#P21-]*2@ 
@BW%JNS3I#ZV0'P!^&.)G5/S8)[NPX]MT@5-;_*<T :$ 
@6@('%UZADLA-=#W7B/](T^V]=1A<B+^4[EV 8 QS]#\ 
@>QDVBP;<:!8+<.-JJO]',896J%/N*VB.U:7O1+PCZRT 
@YAIY.\5;.D"_",L%TK]0T/HFS+;^A2JWC<*PFURMPB  
@HH971ZY6Z+AA>@BZI U=HS\4M^D%"?$*=2ZK\I)#S"L 
@I<F)&-R'7GJZE,B#HF-(-K6^UF<Q2;F_*)L[ON3K?"P 
@["!%Y$^N]08;>^1_LNA3BGMX,Z9,"N)@9Z.ZR'*X*KX 
@NTAY#BX2JA=UX-W*2T1\4*PW :$#WWV:PQPC,@'C!U< 
@HBN!#I5_W:ZW3B\#^N/#3J])(^\K?+@$2' +M533(F8 
@U?- +$!O3%Y:%6N&DJ38;;4M(V%!A#3DX_"MF;V /KH 
@8O!!QR>-G56D#[<-_V5I66+AIL;V&\9#7VX=4H/_QPP 
@MC6YFT)L[B3Z%%BG*DB ^5'&Q-'O.=U6MKZ@,^S$ :H 
@ ZZC: .M/ JXZ?=TYC A<IFW9S+\>@, =\W$T=%UL38 
@)L:$CL01BU5O^X6>V;DK$)ELXP[@[%I4_FMZ 2<>-T\ 
@P"34=^H_=&9B7]#,#*LEGM N"!:$995D@!-^C,^4S40 
@/Y_*(5>"NZTIJD3A0 LW@]^Z>ZJ?$N]I\[8R%07(1<X 
@R9K$9+*9+UL5JL'NQO!SH0N^ $:\&_JK6JO)=(AU(@X 
@1<Z$LPH-4],R?WJLZ%Z'-: 6 J<F>W=^5IIY'I!<I<H 
@2+!-B$B1RL8&"4(WEI'6#R?/RGO9O[B3^_T3&_N5#UX 
@TG"6^1:&JS14=#M\D6KYJ3SK_HM,C-E:K<2+^@F'"UL 
@C"I_G''08S,MN$:,_ DB\#,3<<%/_"MGZ<^1\;]2=O( 
@1ML/+-U_6@'Z7$=J"Z]H?ZMV2-'5L;"JAX2;>B%>Z%@ 
@_^]N-++'O]E)8CZFQ7^K#F&F4P_F]G]JU8R*@P!;-RP 
@S5TPC]WC^4GWUW6R)1PY*$"1E\%6X'%P@VC_%CL-M\( 
@!FQ"JU\^CE&QZ]H1%*"36#%+K#6M;6$) T50>5>MJO8 
@49!-$^7K=7 LAWG\M) Q?;&$T,<T<W\LGU1)*>37?W\ 
@UFJKD$;FK1@&+CM9KE<L%,S;J1V>:M.#)%VK*;.V#GP 
@$UABLS#]$(@#T+'@?0299#)JF+V-UZ5;RW^A[0SP(6< 
@!6F1\+YH_H?Z'$23K3&C(Y<T^)W_'95]*PD1V_^5/Y0 
@G4,7'G-<-+JA)')*6!@BA$R%EGPY?E8#,AC24F&4+#@ 
@EIX)EE[P:U3CPII[_GTZF^W9N5"Z#KZ%.4&_H?>::"0 
@4:\$5.K0%V'(6$$:M'\Q::U8? ]&*X,7B^R%+4TK%3D 
@RV9K;QIP\EEBP>Q2(O]A].@GJG7O'[ND/9 .1[!\[!@ 
@(FITY5LS<S(6I=M:)!$+EI,]1JI>%=*'M\"I[W4 G>$ 
@B/"B\)?J=)6;_U/:C-E$,WRR29R?\DO:!_3N,,25"P8 
@2!.=-.I>M) M$AU[!*N= -CBE,74>+H6A3+I0:0W"WT 
@)/Y87'%US</-U&M-J\:Z**DO,.GK&.22NV"PF_^WZ50 
@+*PBV+ N*\^G.LL;A>>J/J.4&T;RKXVH@1<<6JR\Z0< 
@*Q50]Q)RI!7<0*,*O^6[S.$46#3US9'$_R!VA>>C]7( 
@W5MIW)K2G, O*6V]6YYQ9QP(VKIQ?TK.R'&S[5A5E$  
@0MMS8Y&<X.K4S%&%+L>S@.:=1>3 !8*9?Y33;OMW-6T 
@ -U5?PQ0U"M*93]. @.PLY.@HO@@N."B4K/M\K.RW*X 
@1T_O0F^'I*P%Y?G'S2;71"%OD>KZUHHU>1NC-6$<CF@ 
@X)[& ;!;8VPHLP=X(X$0[:I+G$ .=JEENMT_X93  E< 
@(YU2?U1'W+AJC2B0)2S&>/-)>P;DP,9E<F^^[:F@H<X 
@V+<;^3EUY3SE(-&96+A?OYL:GUM>M//-5P15^/_0Z2\ 
@@.@,I5'>?,(657OH;F."4[5TN$>&]\USU7W!SV (Z;8 
@>WY9: ]A]Q;&U/;8VT 5*GU->7CVOAF_:YZ=Z1QM/$L 
@QM#_7HIV%I2>QPM$N=2ULW% 3O/B'*GU]T.1PXSUL'X 
@?\]PG=4RH:;D1F[4F?'$I22(PKGVOR$SW*WL9X5J^-, 
@JWUS;L1%&1:->3&GN3O\A"1(3'_\W;I=>2K:8Q[#O58 
@?!S-;%+U!$&_&80(8M,<[WP<#$PO(RH(F4&3M8A9U", 
@@::N2T,KEEAQW.<'(.EIUPBS=3N Y4#T]#E:PZ&)2WL 
@*^M\N6#=KUM4[\B-GUW^&=D7F 8^DSIDYPED3 !=#:< 
@D!YG&+WJQ%#NS8\_3*>D>&#]+Y.Q*H(0I4+7OO-8C X 
@GKR'K 11@F]E3B$_+66&AK/1EZA96@#I.$6?N0GW*7, 
@^=H5O +DIJYP?0475 :>37P:;5LB&8_ZUC2VPF>=V1  
@L1-[A=RDHW*@<<Z\_X.X4EIQX0[N$%8]8X3-P/[,=V\ 
@%UYHZI0XC5V<M4);B2\GY<SN"#-',V050=:2*H1+XJD 
@M= /D@DXENJJ,B0]XU+?KWG_T<UI;!/ I@!P)XK9><$ 
@:B=@CDJ\.<ZEE/H\KN(TOPTEK- P@&V\UL(Q] >'W%X 
@.5+Q@G+8%=3S8O@+XJ(2QN@"LGANE:C"X.4TM24+6LT 
@[A.7+K??7]KW]M>X5_-F1[ZXC_<S9)?O9"+D]?\PNX, 
@'7C4.[341O8[7EXRUWA^R=5%(3CNR2FBZ[*#M:Y^V\4 
@=4LC*'WT-,*8V=3DJUF%M$V1<L;;UHS;&_.)*<%?J$P 
@#E^3,U+;J*F^Y!C1UKTV'L84;;*@+.E9*Y[6?PBL-_$ 
@Z\PD"U_!PMF#:FV&ZK(PPJ+=\63.<DOG&Q]GJTD;9\  
@7(N%JI9^^B;EC6=N/&B_1Q9ZIA5D%Y';UNM).LHM $P 
@.M,908P!2GV=9->_>8B=@GBSM?R'2N4]72D,F89'1E@ 
@K:PVM"*[XDNCPY[OC:1\DW#'>EW;_<2-1T1?V@@M(ZT 
@M^B= , 1FHFE%.Y%FH#T_Y3>6QL,VA/Y:/PVHOFMLC( 
@>T2Y]FD\3/MG.Q;SR3_U%(E(_H$B<%LUD $_JR=P6\X 
@PM@:*>;LDA,)]2/.+%VV"&S3QS1.E":VA\F8B]"#,.8 
@X)<;['219"Y:D8848EQ IS7"D::ARL__-&F3L\,XS.D 
@DA?SX"VD,[K;I.3;6%\7^I IC*:<4ONBPK3<;K'<0M0 
@HG)47<,?3".%@\8O6Q%V6'V.ND9!<<&IZB6FF%M"E<, 
@U%XF>O3\H,9, 3*RX@?6T6!7=PV$.&_)-..JU32*+ST 
@]"HXNX*6Y4Q$!7_3T")8TN<*RQ1'#ZI%&'6]78JEG]< 
@*W7'EQ,77JKIQ4WNN\6V L^_ 14G:PT3A],8:*QXB"4 
@98)NSH(56_):IL_7."V2QGE$,.&@8D'7^3&BE?-1+^< 
@:O>B/L:9BM<$N%X0_,:2UXX):X?!AC_(Q&,IS%85(GD 
@4Q@O5Y]=D&J+$KNYB8KP;XS3=%QN;9A\.[10;OETWFX 
@L\TB7))I.Q<12^O5YI]3C?$I>0?5J_8P7PL;^K]8['( 
@-E37& Y>GL>M.$L(42#!?MFJ?68Z7;-XZP9A6/DB6)( 
@>J1#57%?8S!5]T'K+^2UE34\2WP(4+SZB$T%M6_DO04 
@;8EUB?/A 3V[KWOVU1[R2OY+'H*S5M'()7^X)J=)[;H 
@XSQQDS"&/0J[>TZ^T;4&\_^*42^YI;W\*NH'].NRUA8 
@4?H;HTMZ/#++Q(W0#WYS*F2[*7-$B#(Y)9ZS(Z%CH_  
@=:2>7#5 [[Z'4VEW1SSOA%W\"\>K68"'G;E>;1$Y'=( 
0\7F7M9KZB%L,Q.)%YSHG;0  
`pragma protect end_protected
