// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HI\ZN7MI7;3S+D;1!^3_S<(9HO#75(SUK8(DB-$P_AW<8SM/_> PTC@  
HIH4JY2UT Y@^NAO<0Q7CQNLT-3Y:-PU'N-4*I2IG)$@]_%1.7'F.H@  
H,J8Z6%!M,HV0\!+H1_-L!>OK3+75?=M)32B%0=)",'J@7<^)TY.9X@  
HX'9\U#RFQ*B,75L2YE@7; 6)9H-IF]@-JT/+D'6&BY&B30>]^5"\?P  
H^[+2-[H7#".N7[\<IJ2-F%7'*+Q/P4;OF<:FBH:_/8I\ Q0*U,-' @  
`pragma protect encoding=(enctype="uuencode",bytes=4464        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@E7%=N<7YW@>]09%ZRF6CP#\?S#X-,1Q)LXP'B>DH/:X 
@FFF J9;IA@ '?&TN= <>FZ'4MX4@G6L1I#@)VV:?5UD 
@O)72[6_,6V+9C&8:6DQZ-+'@$B!@?P;MHS4^W[K&#1$ 
@^4!CC'G1+@R]A,3!)1ZG?GO?X5VOQBF1#U;DEX8NQS8 
@F]RK(5MZ?-0J==Y!G]BE72("YZI9_!I(*I%B])V=]"0 
@=V]L\C6Y,?^CM]G&/H!;*_T<%H4DFU,?1(2UZS&)"Y4 
@*?I'.L[<''8[U+_6Q==ND(6ZKC!_%D0F\LMFCOK%8Q, 
@YJ?72N!-'U-_YNPB>#:367]868BR.J@:39SF54:9%6( 
@]-5^\TE,VMPW9"Y17&LNR6#ND?\69)ZT>71-:YH_J)4 
@)ZEW]6#1LNZKF*4!G6HY3B+5C,E-N &-$A5*J06Q7S0 
@1,T._S%K%("*)FUM"HCG1?U_L8(]%U)M2>02)[X4%<( 
@:(N:'EKD-TE&_P0-*/JC-J43,-\0))"BG]=N!5LJQX( 
@%GCZ/TAY66IAYT3'*'HN4'!:FSL&BFL?B-*1,S34$ML 
@_C9VE$-_V0I#TG%ML?2/[O&QMD [?NN/MD1LP/#JWX$ 
@71!37)PC-S1UF H"!XI[C:A.)UG%\#C/&]$PPKVE15( 
@:[!=6_:.G@B;N?BD=AQ<2\7&7.4&,)!89AY:2=5EKD\ 
@16QJ8W.M R"Y"KY0I.*ZJ=GF8&M;28BGT@J4:SSM%X< 
@E,S=^Q)PM3I=C'/[T;7&9?0[]P;N=871C2X+P^W<,X0 
@S%YG7QDC'=HDU2'6G8[EU:^TNTXG-L]IPMO+U]MK'ZP 
@N4*$7@^6H6_W]%5^,%0*H=91\&3>W(*95@X*&:V2G6, 
@&MNA)L[<E-4)/T1DQ^EQ[LW[/:EGG>K6N@F:6*X]"Y4 
@BQ,GX\*I-J>!0996_#.46+5KJ\?;!MNS_LW'.;&;)8< 
@<*)C^ROB)9G]O^]!KP(M,4L N]J>]"4*%%415:2JHLL 
@OINA)99[P1EJ"4@HH %80^R8(J'>P[AB^41(F76:*#T 
@S_E7C++'2OUHT68I\+F]VMN#M[.;VT%)9ZJ@1-0 J*X 
@D+$<C3CG-KDA6S6&5RJMT=U:MC00.BH3+W4L:%JOKZL 
@_J]Y1TZKQ4U*[L,[6EW@X]K^Z&17[  :0Z."IAS^4J, 
@J8!R,%P2X,E. JR/<WH5.^UDL&2J%Z@SM,WCF.[$C6L 
@;4>0P VPH7_.-IMSQBMIO*IJ$%TF?AQ9/$H/9C0RXUX 
@2*YL:#<=$,AL?_].9_(<20.O0'AO2!H<\IGXB=:4O@L 
@<'GL!.1N;^_LN):43*O(DZ&8TM6Z70&GW9YWIXG7\78 
@WF$9WN=;'O12<CX0NM,?R.02?:T\_Z(9 JU#CY0!F>8 
@-]AG9+TXXG23%!*\FI*:4J$)]!>@&A)^+\>,N=SG&_8 
@$=<F:B9.*6=WZ.I[F9WR>PX[D<N6S=M]JP._6 &JJ+H 
@.]?>9P/Y&$(<QR26@KSVUSWC3AML;+,C"3K%DP8"]G0 
@_M(B6RY0E]7:%L7.@EY5<)<S8%;W#&!>N[9#S)I10<< 
@8W0/;_]9Z.NK^T7"R)6THS-3-%%'U<I^:<6QAV2M5+< 
@OV2Y!_AQ-%= ).\-K:9]V=IG):"<87;W+\B%):-V+K, 
@X:WY1_GIXOP$XNB"(<4A%4<\^'45+0$_X&Z*0!!=RU@ 
@US_ Z5RZ=7R#IR1O +D=-R8-Z1\SUD&\$7/ ,@W>LJ( 
@ZKX/!:F$_S1W2X;QA;)/$?^"=H9].1Z&SU+/*-]+!S0 
@:#Z]D,U&<BG>1 <:TM4I\W:!2/X1\+*PAA[]6)JRMO8 
@(G<VS;TA$UV=UJ:YG?-0M_[!-K>?[$?@\[3LX0Z"'.( 
@E)S:AV*@11"*#/<K6>^V_ZE9K[XJNAB_\N, R.[9>,P 
@2VU+&#E,1"AXH$:*ZNE\(_^--91)K @[83E,O7K%0N, 
@S,"/_I 7R%CO;Y%HV$\N1%GSU0$^XH]4N2W2$+7R!<L 
@(D!V[ M=2IC;,%1B!]B:EZ;.K_>50C_?K)42(W8@/LP 
@I$$_*&H3>/?^0@B \+ZB&<O^G V-G^96ECJ1^2>(<!D 
@39U,5028C(TEA_J"XBT:\3$IOH^'X/?$LH!*RS2Y/<$ 
@G]SK05'] M::&,I(0;:HL<-^_TY%L".KRF)9-.=K^#P 
@9-[X-6:B5\R*UYIY[9CN=6NU%<<1EGF&@Z',M1!+C<0 
@)090+KI()&933T,Z;T$3P"7GJ+^.$SR>D@$6QT:A:]D 
@HY/GB2\:3'-%/U/ASO5X,8_ /N;-M0@Y^>_?")/>J9@ 
@LKFR;)3D\5:&W,A J7PP #W_ +4DBS+_?E3:LL8(^-$ 
@A4J&15^8RVK2)Q&7$D"%965J;T4,R44<=-[>[ZL#5_D 
@M9+#G[ @Q$]S-AE1SR&9.719)%B+U&UYEZ#D&^X2>YT 
@K/8R'+&OJ=$W* N,YR/_)H9"T!'RVM;09R! 4?(FIVX 
@H?7+*#W;&?CM!)3B?!'W^?(W[T5B02IQ=R8[AI*E]3@ 
@L0#@)WF1\9A(-L<$[4?6H*:N=*_%3=R)ZZ.#2;Q>"I$ 
@2YP>C4$8E'FX#1 8,$RR'3]48\A,PP,:_S!1[- U#H@ 
@\905G1]*4-N) @KMZ.S('4:]U_,H.^E]P(5SQMPPR^4 
@27.H$83/#/GI(10Y"O^=U?705I (_P+%OBN=FXEEI\X 
@=!K?02@1-*QJQ)FT6Y9]:$ \DYT-KV5Q0-'+_#8#W]( 
@MK+98A'MRO)I,C55K5\&TGF>G)8$ND:-'""PNR>&E5H 
@55S"=BJ4\%5\ZNQVK%&.G]F8J,VSI[J#1M:TTB/]D6( 
@HI)#:,DR"K)"*O6U:S0 .'5'[[]T_A#FR#[*G.>_BMD 
@]M36W)F%=H8OTW"@ 8MQ)92@G>,^_V.E-F15=*-8!28 
@D3F8[IFYYN6X*P>UN+UY/_&1V0*_WQH M<"HMI$FP!< 
@VX24O6/XJ_?=D()4NA2X0/B;>(P7H014EW+W6W=Y;;\ 
@+0^C4IV0M*G1SJQNG(I[):]P7(:_2 VS&M4QZ%?4EU  
@F#T&H0D*S#M\<N.*T:@-BGV1:4]OLC!B.^JK'839+70 
@.\>?Y W<*[G""?"EH'=75W>9(%\9^$K2:P0S7<.J1@D 
@0 K>M5EY.F67S;CV8BZP"[S,Z"!PP.WFQE^8<X_E&"8 
@Z[".IED^6EC7QH#&LB5P%(XRJ70?Y3# DQ(7L#/SU2( 
@V>D3[8[+GZPEL[2Z8:(ZY&[1=WP9Y5_KG0S*M3H?,#4 
@V1+4&8%TE%;][P#.C1I^68,:D^UK70I"!Q]L^+VJ7MH 
@XC_P5X ZH^KY'F(T]=)=K1DV4(&3#$"6#"4#"<R<YP8 
@M<LZ](J^;!2;?GQU)4"G3&\-EP;M_SN00J60X'[ LU0 
@26TXJC$JMIH$(ZH26$GD&Z) ^89$#?"!(:XG0%X^PI< 
@RH'ZLTK=@C:5?/L 'I_X-[#%FZ[^_3(4:[A'?WX&#1\ 
@-:T?^L$.0O6;"V$D"(K4<QF@<CF=*JX7G V5<MY"ABP 
@PP=JI:30H4E&+]5:<JW%MO],B,-#$D)-^U=;0&03^9< 
@/'F+++/61[[(8,_I_A]Q^W-==1JI\K6N8:I"_/H1:P$ 
@;V'N:858 =O%5PUW!X2WH'_^#[>-ZUR@'=2V3*/X#WT 
@+@]M.6BD:7CMCZB$=JN@ ^!?HZ%'H 7+4)K[*)O/$;T 
@E$;M*5_.HH<)RDZMWSK3BHZ1\*B;]-V*=7U@/0P!G]$ 
@][>/C$LTK:9S;:D/,=F3<CD48;O&6L#'T) /TC5H_X@ 
@ BW39D8,#F4,6)5RRQ&"'JC.K.E-;LD$2&7'F#N(@NH 
@#3' 8,QOP'$FU:1OG<P="A?AKR',R,S\U5(#HE:M:TD 
@]1P A+"'42T(Q'6N2U?<U*?C6O?WNW_ ,,W3_D\B%MH 
@.#-E[/4MN:XK/ RVJ&XXS;%<E_)<IP_HG:=KFBR3B9P 
@8;")[1!B :C[=^?+WPRIB%?^$W,J'VRU]V!, (Y R;@ 
@(L(HO5LP65@[SZ)=,P=&$*DPV7)LM3G)Q\%2IF[=M.$ 
@7?T8^DOL#8/[J_S<L9*O-MO+]H$-AC-*O;QV?,&*-%$ 
@@K!QYD_MB&TF>0)AL])2O-UB1S\"<75"A?QZU6]6>"@ 
@U3.J)'1)*[R'KW14HO248]M\>B;>UPOJ4M^JS<&48LP 
@J.46_7!*HNWP2.1(]$17G'LP$/SX"FUQ>!(+X^.;_RP 
@B9X_YNF87,# #8289!-^04&13CL@6SP2 D0<FV7JCM@ 
@4[.RI3:"W%/W?+X[SQ1G>6\D;M1O,;6J3R6HGT3%0QD 
@\;&O/)V,VRRL<Y(1YU6+R&<@ PE6!(UL?SN:=J'!78  
@60K/&ZE^X'=SA1'08[G^,, EPV%T<"O*2^R]N)FV)6< 
@Y%6>&*I-]<X7V9,E+GL_R.OG3\%TFZRXD].+!2O<8G4 
@^ZYA%()C:&R(HE)#T*61,8'EU4+);41.JFN_!&_Z!I0 
@8!TE-9""KG]DPU/G=Y&&HZ,+.N<MO0/( P_4CD!1M54 
@?=T:^/<Z. <B,E@=T1&HGF&7]IG+"D.A"^*@/3H&,0( 
@ZVLB)?7I)6EZSWHMG69F\Y")"M9E;L'--H=9/DNOD", 
@2:Y<EIW9_2XB\4 C#KBR)^EAOB?>]VJ"XK0>@;@%F0\ 
@S..4UK>*KNKF(!-2[IKLV#JY;)0Y37N%Y'0Q7GDY4B@ 
@.A2QOK)KA=I8D8C N'T>,$KK49)"9>Y >K[4]1=B $  
@(+^Z@_G9P^#&A"7^XYYOL_(R770JP,E;7\N6G/$U$NP 
@\A7E6(/*3\M_Y?PHP&Z!](C8Q2ISG?-,)!QDE:E<?/< 
@]E*L FP(^T-4<2"GE33O^$O,IV.UA=SDA,7UU03X$V\ 
@=C.BHXU$2_]?7J?=O1XZG]%)T/O5G"!3Q&#_N.GBU=( 
@1Q?2S]5S8D)OE5E?!FG-T%5_:H19%B'NC/*6Q/F(FX  
@"Z.!'9=4A@YB/^S>PUS]V>^^7Q1N@L>X@P?@;>M\<&H 
@8H^W%(Q)\$WX5SC)+1*D*QYUA4@VEB\W]95U'EXFU\  
@9B1T+V@_-P(A2(-B*IDGH<XHESFKOV] ^!KY$V8U\8, 
@EBOQ<<%E6@<7'?(]X_;_%6\%7_MAQ/ DVQM2O8OUKMP 
@]];D"O'E+F%7I/\B=!^!;\R O-7P9O8D2'$ C?LILQ\ 
@YKK<3SK54,'8>G.:[*MLZ7.GWG;2<*OM@T8FD776ZN@ 
@4Q]-CN28EU.&M81S>SW=P1W-A==9V:#_6=$U0N\++'4 
@R/J:D$@]C/FS9F7[F2OU!3GK2?:W/#)N\N>TEIV#4=  
@&TWWOMB@7;:7PWA1X)#KWY!!BK,_O!YWNY:J8VE[,PH 
@>4Q&ZUS:"E1?BGSKFU<8"_)]ZE^O5DP1$!OKYP1 X*, 
@VA C.L49V%>?O+Z-0;^L5%#I_I'N2)&H^.-+W[/,(P8 
@&H21S-N]ZH,K!/YQLNZ@,M-+2W6,#ETST<IM"3KE'?$ 
@ML(-2\L)-CC9F[59D*E7O)T-PFK1W%P_C*(8\'CI 0P 
@G4,WF3WZI--8IR<A<'#@G*FD%UXE3COWZC8W:G!ER:H 
@*%Q. -W%4K*E ^?G-C;<Q&_(/]EK@;T<EI\T==A=OVP 
@,FH'[0O2Y'Z$AY_"<.Y29TA?:O1\=BE=\7&1?1Z&.&$ 
@:Q<JXFAOXVJK=<>W4!J$;<,V^RZMVOV;Z.DH6[33WDL 
@$_:9OG0WD1J3_Y53ETQEN6+,\\AZZ0#T&&_])III$ZT 
@D+:]D#8B*7/'_J3P@+VEH/!\2&@K;AQ[HBW3NC:1W54 
@>38:&8MHG51UF<U^![/1WE<6\?.CPY2W!-]ZZI& #%X 
@.<90PG&&CQ(2H,L!<Q 3;EY#MW5RW1;!-]7&@198I;0 
@LW]6D2-93/.P&Z9E"V(S43*E"Y./$G 2E9UUP-@;$ZL 
@U7"GIR>1"B../ GT67$L;+F>=#DY4GF?ZE)#G>5/_!X 
@+?<^WO8L*BC@.F#SWJ WK,2P&<9Q4(K?;D#DSWO-8,< 
@&P!!X\@J=MMGM5>:A?-*] \Y^$5[?A$BJ, S;LW>G1@ 
0&AHYJ6+_C5@P]?-JW=ZTLP  
`pragma protect end_protected
