// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:57 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V3SFoAcAV3ohkcyVzpmTI5TWsirz/TlEwUDeKYvhSbbqSouffSyCxLt49vGe6luj
pV2/VrOj+najIn1wCPwvlmU+NqWbqHQGyZTiEQT7e7jIos8WTo/LGaZ+xTd9jAqU
kzhDkSDbUh1yEwp2qCZ+YQK+lDkl7QlhleRBHw4WOGI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5680)
U9xIZWPsBVprGGzE9v2BbshL6OoYcvUIq3Y8OkjGW5C+xwpvWvxduJSs5Bfpteq4
1pYnEYc25OuXj4j00jO0Zmaq8ywVaxllhvRjmkT7vCfw4JgS06uMPGj+/7+Ql+EE
yqxkrVPs8+pOMSycCW5VMk3yj/36F2lI9hXPZqs+MshSbzpgK+t3GNGh7uIJfhw3
0ycTjDEIn/0M9J4LitWSteAn/YI/GPziG2A8Rh1sGMWAEKMI9PJYhzoV6/7K/CoH
YIunAeQNgiluRDurr3nCgB4u+P0MrjZCwZ7KHU8MSD9cMn/HWAB/cY0EXIxbLHrm
leplVsqzGogJiM+c2qZdvgPULaEL5iQg7VemQrrCFToQl1G6WYivDBUaZgcJPZiP
yC5Qv9j8EOIrePnyTXglJxwTVjE4C06DsMRYmzy+lHm8TlrSj0FrzoHcdkA32QSl
qXbPznjD9qv2yJXWI1lg0QiPQW/uA8M/QqLPRQjws32B7aUqYzrzvMfQ/PTfx/BP
Sf4bpmFHf0qOyESoMWfi0Fo+FhGOeYqG74RCcYENImmsBjxYTwdIUdg/5vSfMzOC
qrt72QIeIqyfDZ6VfKg7QIvk6vuZtk2BpSRn/+Py8wmopfcSlXJSCdoS0fgO2nnn
QGDxD8x8l9/XSu1ZoQ69f6UTkg+U70c81IlbqChBaoegBFvCieSqDUKAFVPMZXdA
je8Yco4O3vhNIdpA9KC7r0Lmw07RiV/JBhzoE0Ct1P2Ra/02t2jLdeh/qqIS7Cr4
Oflv3RlTFHfM8mB13w4bHMSwQ8/JHL7+BYqJDLd11JYAh62GQzbhzYsL+2WcnFHn
t66GDX7trLzNPwjNMBAu+5A6rXNGsRk7D5/a34JlW8SQuub+yvBjPkbQ0EQmitxP
eo7219xe7WyqdIdqs6+Dqq0GmGHIWf/64kzdQwqrHre1aAydrtJDmHBwZX38sql2
hfGvaWJCqR5sNU8E9rAITusubh3dAjr14mHFdk/GqYjwxrApCmZDQgLOGshT54wl
TEreTjm+PPYr31s0ViOcSQf3ucLQQwk88brZ9aL7u3NH5GjfdFQvxTV996P3mVlv
CRaKDsE6Do8GwB3aOQIdnQO5kleltskmxeCX4ZNwe9zaFBIzjPNLLowuK5FSGilF
bF4+E57XGxuJdVLVQAgbv/UCqqs0UPNP9yGMJVOIcYmGs7xX8oDO3kHU/iSIiFF5
HR6hi4eT+LKjoBetDXaDDLKc+B8H8q0axpNFwUmAzKiBp3SegA5siFzE/b9pBZOp
CJiUbKDv5fsHOfHZFoOWF7kF9c4J2qI5pIs88M2HykrXyIW1XbifVRvXgj1drOht
9GSKtKuJ7hef0y6mt1VBik+3JJL5PMJJudYEzjEJY+tRSIp6q6KG45iL1KZElMUq
XTNFRrf8kYNchnOqZLoizIgRdLsv1LcMZPto82F0E47B/+IW5wRMJRy0r3ioL1zl
GKPuVQg187IUtYv32CAHtOe0rqHRAyQzlqI/EGMiKUL9hgIN5l33VsW2L3hgCIOf
uFAdpM2kFrSRVYUOkjj7Mv5fG2m5ABTvezDHweRb7WDblAeuzTpkhx+9HxMXtqja
bVcqaAyRst/B1nW8O1gTVaE6dDJKXnTo4L+RxFyM4gDtAJ1YCf/BIxhpK7ZKSbMl
OXAe3yPcxcWnGuiEfACOhjvRaJVrNe4l1YY03+Rs5PHmwKZXcARLho42rFUvJRkH
/lFok9kQ6Dr6WdILjrmar8llHehfKICu3rrNOEwowXObD5SYC7p9NQMP1agRh8ot
8PsJPvUO2X9GEz7ZNAC+fL4f3K9kcw5dP0jeogvfdH4pct0nC0Q8Ap3cWNhWHh2O
oALYGDX2CzglxuQv9OkEClwdV1Nzg+jUxAbkOArH4nhW3QmutVdsQ7OQdFnrD19S
i4CqXxsal0vNvAPdzmL6qXCFOtx5Mi/NvH6xafhIRlwKQTmYmBB97jKtaJOFls/I
UorEmNJjPNPwIdGeUC6h2N1/XUAWZ7YroyB62dmFwwOf0jk1thdXD/89k8bUdPi5
+Pt03WNWz/m4YRcHeskS0uA00qrUUudc3LS9O0/D6woxZQmM5msHLB+kli/BLFp5
kK8d0Io57dtMBKmq4Y97FdyW8N9f/BlKwc3eMKdiVBoG/bPAtUebIzGE1w6rJ1we
aD9ht/m2x5Pxz2wrvRVkuqPbcpE6xf+vh2ljchpvyIyjZhCECzafHE2vA73kwwYJ
256XkZ8GeFqkTSSDDVmUu2ZZ66sj769h34GP0EXzdZjhVfZFHt8lmqLgBR8b73i0
lQCm3eVMBdK1PK8pNe74Zs+7P6jdLLH55M4TT2TcK2MKbi3YT6cEafDBOxJfooOL
DsUagx1dIovv5hKXydJHSD7K3NaLE4qKKw2nnwGxTPMw7MqepBdgtB9uW3c9edrE
/MugS1bRTeEWjvgulQ36FKbs5/C8nvgfd89sIIB+dUa3xtE/GibuYZLpwOd4/ij5
jDQwnbDRQATV8OD9IFLsucKtAxunpRXitSu818AcAorhL4PYo8wEq5ep4C2A11cG
wlxAJZ5NqjLzmkwpltaa0fsPgTKDRfPzzil89Z4PdxDc/b/67uW2sgCh/CmE0jFs
H9CTRy3FU1C2ChYRiGh2XMB4n8U+HDZf61J5347q+ijk4Lms4LpurVBsg5S9aiHL
hA9UNsXurVrQqcOm/m4xPAsv6IDje0NWRfi4RJ2oWS3SR3QI3t/wRCnPYVQi+F6D
hdA8oNgev5zpOAhZzDTwnHFLlgbtE1dgVEGAFeO4p4YLQhFs9z8otnRWjanvOcGO
4nj/mFCrZrCOvFE7b5C/qutN6UTWYru5C/JAFaNFozxgknBAQV2ru/zqS1q/iJP6
gr/ioX8qD1dUpuLYNg+vo5xX00eOay5xXmX0l7WcfHE9PSe4uuQFj/SnqIygzJU0
U92IcRLwjuGlYVq4kdw6AxnPj5VcyFv7i5iSQRQe3Bia+OSsoO9ic6bO+192VatY
ztZZSJ0J/JOCRsdLe6Tpni6fm8rBPgh78FdDCjKRcvgT13LBP8CA7mUCjFLFOiiu
sq18/YkD2jRuNnhIKxlUOTzfQh50zhKd5/LNvq2gfFieK/2BZI6Wpql/AoyFs+9/
Kfs0kEqKgrXelyW/E6i7vUREImobUbLBLpUmPDe962Ni7PP/8N+nxMzcCXPKNPri
8QN868DBA4ldjwary0iLrM0UrdqURe78u5ZynZFML4EjAeShpI5uTnBg7t0Zmrpw
SjXE807Up+F25J8OGVB90HVa0mSQxSvAM8WaMjfmGt+aWh7DEQaas0NZ9T1oow/v
3EXeMvm8X/XiV5kInnz8hIJMBxVd6Zvo7ojoVDco16D81PYTixTXasqzPPYY3nzK
0ISlgGH3tBLb7ybDW95DhnsHh291Cv20h0XB7+EpZz2x2ChZRp5eBONR6WNlpHzx
TJxd69ELKx/A6MyEazuWtQL9mkYt4OeEC+oAAbE0ISH4CIp8X3MxeNA3o3vQg2Or
PiaE0Tv1lB36l3TTQHxxxiElhavchUEGQlm1UQ+GFJitZC8py5AMGBzzqFHBlOqo
C6sBl6+s63/hVmaj0SRpDNu1jBbpnUjJsLEofBfme8Oz24iZNLo7bV+0ywTwWYyp
PnWgYv6pRT7Syyq5+CGrP8uXb/n8j9IcUQJcPiiSzT0WQJhIQvvTnGx5p8VlE6xY
Aw4EJey2DV5gMFJWjDzWHZamLDe903pPFCpekTPgdaMD+oSGcInIFlo79uoTcXik
XYwXNqQzKpdSJnO7o8DjSS8Q+sRqeK7NnR8a4FPhn9O0hBT4svwROvsRIY+FXmZP
5sgE8HKUzlEUHbK84a3aLeXHOjOpZPigesBfmVym+LVOynz2XoJAiEJJooEUwwk1
KQH5Ct9zK06JzxBRfinYU0QFjK+8Fg7HHJuMnTp8T8+1ADAEYADofHXt4jYAF3yR
vJh+As5CiryvpEEHwrZFgh/f+9SDuFWYO7wglggLAZKQhR4L0KIxSuPrwT0hWXn5
HNczekBRLMJKoONV/xLGo2a4LNByqfcYaXQ0k7jxuXZ7j26FCQiluXDzvjK5EBoj
eUHb/0q9OujdbC6Ehkgg/VHJ4KbDAwzjqg7Thuv6fuBcxcSNY2X03MAGLm8a7+7q
biICzt3wXbArQieoxD27330W9w1Z6uKfJXmC5hxd93XHAcU8LvjXJWLnpdjZMXRW
+iDWsd14GyxAF7XSuSQLtDTJI2wgbAnGMAzIAN7YM7UC8SIGtf2+wbEEIjyzU3k5
buSGN0iHX01l0SaiwFNgDlb4lj4CGHR+VaO92F+/8zOvVaTtiYYuTAZSIt1qLuzg
O19aLQzWwx3v10gZ2zS9LBJwxrQ0SCZEUNXyb4zaOyjJnxnoa+qTn1H8cHZtb/Ut
x97nzo3i1Y8KG6NePZT+cYpHD2lqxLJoWY3tLWaYrr76pT+CkpHuW7xim6P93Z9z
5IQdG1X/vWAH9O33aotP95Ub5wSu9omla8kaBOeXGFarDcbr3LO6AxLhhBtEnxSz
tQ3vV7V+vQRFXIby5HBGH3aklUJhfWtQScq245+27kdcNneV89rRkQMxIrzk0FZn
LRlTAQSU3MgCVOO3VX2ssnla0046Bl71xLNsgQDRSh4N168Ze+RtNjyfU7taKM4m
udGD9wjTtbotWZfvUSNvfNE4P8IAaqdAyYccJuKc4ODvmM46gHSbWFUGsL/QinJy
jqjK96MyLuhBH1RXcr09x8AFF0iB3vm59bFSjBRKa6gm1rt/Y7rGSsgX343X01u7
XHHbiCimce0ths8pk/dv6xtZC7Lq++sKgbm1uScT4DJHQN/1pSHUjUZxuzmlgKm+
wsT4q/3s3N5bfdl+vpYwnTtz2ijr4sUTbYl8pfFdqZq8hH9XQ6TlnrfKGFk3oJlf
Al7vcGGvSag0t4LY+KwX6iRMwbNE9gk3wpbAli3KeIIwDqbI+KFUGyqb5xGpfYQO
i5/oO3iAe9oilowHNJtZPJGHxgA2ZaNHfz0+PYYfFDqx4K6N2DheVIETP3ezomuH
THT5pfnw2DJUzQEkW7XJMON9sS7F7l+a0SkrXYBtguhUe/It9N9Gru6md0ct7esK
i5BaYgDuIzxY9baheoRHAsgwLDkcGz7kZ7HeA8agwkwLWzn09NCI3KEUbKkeWozq
a6U9ikrdL8jr+2fGr//uqhbI3ZZkBU4feBecuwmot7B/m6ysHycDNaHE28bs7+J7
UQ09P0Gfb9Ml3rvBYmG2A4gonX8Y2Auv99z+/2kOUA/rf2STLwNQei4AU/PYC/Xx
XVUtUJ4wfHn7IA3t5nj3eT01RiHUbPa7ugfzH2jn2c/rVHP1BIixbsmhwd3JbTE4
EeMOuz5G7cgwfBKAE52JPI/uMu449VZvyRpZ4Tl38EgR6gkRgpCdbWfIYfNdO5gW
Qhs8nGiYuMOQ2P3RYFt6QXs4AzPqof81JwM5S1TvDKwwDiwia6LbyWHudj5J/Xf8
vkkeUx9AwSErKLffC91G4QGLxouOBc2wevp9IFt+4UJCA/aI/FpBL3XxOG9GkEoK
z2p+JkxGf+oURakkH9m/KbXi4xiLIH9R1XQC7zKQWdjAizuIfbyzV08xmzX0KqLq
FJw4vT7Vzw2F6Wgr/C9ELAtC+p/2M/RfoKeDf0oUIZLQcBVrCubApMTsi4zh2V5J
rol8/Tzyw3f3JR/YXvL6f/4oP5EaAfxyFI+T1z87H+9z5BobmmpvGbx79VN5Hfvc
BHtvRDcBIBrdAWVlax++L2qPpMGeUk2ZvR/a6kCFaiat1tV8yVmp4WXvYtHMA8cy
TtIyhsXa0qlmxYHpFakCjZApwETI1lzAk4rP+hcIZY/yrrK7TeyITosiuRSlPsDF
xjWR3nsE17ZN5a8z7px1bEIsL0ceqHjo5J9VzvNl7nWXz+6qSBOnk+Ou29EuvwyP
U/aAMA9T9uooO5JNvn4QGule179la9dG+MerWdm0qO43kJJLdjclwRT8GH0Oflux
t9CrXIXtTG+bwz1ASVZnNfMCxm0n/lMnC3GpoOhMJtotJ9AW8a5uU3J4sHwxRFGI
9TcfCJhC/gnTRvZJguqHLS6O79MghyLVDWO4qlIi7lG8WmPKBQcmnltIJviVj+NE
o7DAdF4yKq2MKDlzfy3j+NPzAVi9XIz0P12bQqES2pyAG7yqGqowTldL9nJcUERp
ERKwV8a3ExulVJIlK1hhzCYG6ndloFhGdG34a9a3e864yyAV4hk8WGUfsHJNQ78c
hEv37EtZ/+dpV6KPq7PeYuKIOLlFHpqT4vLH76VAcJI+f1ufbi9V3chI33El+VLQ
95yXkhRa6D9m8Pe+AUmiCp29AD0Nzei/Ano2qfuYJzBKPUMrsQgihcgKXXjtcY2y
5UiFcIRPJGjVBKQ6sIOCFHquabEm70bdEG1uDuo0HRO8CYwjsvIX+1L//zykVXhx
ZPci2jpbXTYP2/Hh8wXt8B1dbBno8pNHksjGg4XcCWW6Q8VhbjHoJskEYKLuDjHs
zaa2ld3Z6dQ6evlO7uf6u/Hz283wizw9O1AoSFKlPpBTko243ncMhOEQYgrlijME
Qmfm6YOH142UyhOMnPZiysjzTPmgaFhBbjKLOQzgJwTRXdQb/Pxkk0cKYPaLU0J0
2ZIlA848FqX/VxqCrXnem2J6ry70MiP17PaUupZs7JOCut1nqTvFNyFcALs/Rrjw
hpBZpzVFBUtOvF9epAvLJBwGoGNIiNF85hBwJnVqjVHDPS1cpyiQ7SU7x+Svsmoe
8SuhPryh831QXU+Ywdevg0ozxSpnzsEWmVY8WxfAEpgh4gc4quajYkvcJAwemQlh
2RHZdPMG6zRRh+V7VJaDQVfgTC3B7gQf/xpqEDzC5guMIzXKxAA9qTXGESnm8Xdz
RWezfv58B73I/iiFsxxi8cXECxO8pcXDs/bT/4kl7XeAp8xrfnFSrK4I6oISTQYM
AEYx9aWyjOE+KnEYqIkZD/qUF1C2X8haMXC0PtpVmdocpAgqYRXGYkSCoqLp+Ozu
drgjWrGdeP0yXI70g+2tsGuDCKQsTRTTurknT9WB1E9OBpnCljTx8FBWda6lFpVB
CpR6hxR7L2I72OaRmmwIFWEMd/xmfFv0VdFSoEdlvffnmdkvBaUrddeDfdYwKIOQ
gl4Xt6NbIWwwq+g+Nm/aHlPbphefxPd7F8xmwdSqj+1U53P+J/Jix1d8JnU+DeCE
wNhOUAm7A/qXDTqTYZjXF3+LG5HFTnilrTJ8dGR8ST7lADb80W1t3UUDpzAxD5Jo
6tI5pw6J/Va1OzM60y5jZ+fQquCGHaSh9W58u0oQWNkG1BhLKEZtPjQ54jLRgCgB
2X+Um0dhiEG+WmL1ZRJ/RBxXraVdk+1n8WfM1ohf6AG7g4/o5loclAX0g7Z8iUu9
slWGYkvilbAf6vErGrq7iWxBc6kDpqI18OhCOmgewvQDrmCNLnpI7eU40/kzEjJX
zsBdmr++B4B4EiXwn+zMcUF1sVSdi0sR+QQyoJrtnWsXBqzcbFlpuaSq/SfhXkwq
DhcsS0RXvq4OK+7aVQZyKg==
`pragma protect end_protected
