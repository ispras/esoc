// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1QOKAB1LXj4n0wX6W8Lh2f+6PJ+uHfNDBmUTTn5huX8wxYZBlVdadx+nMROqD3dHUPrAqj8doCOm
HNmyZ2xuC31LXm8prC8wcr0nRVJ42+JrgRLbw4/09VcAw50tn+VKg5rAC7kVOCLWICjofQWiO1hq
4HwP1k6kMCtcYXyDMuEcOqFNGwbu2tptyNSrKwIy7bYkGk01oq9ah6P5/lwVZJl84fWXiJcFVaij
FKzF8SvnMvUAipa4Y75c/9fVz4308WfLsFqchw0bEHFU/YYMZwkgux534AYqjKyLuPNq+G9MIYF4
La0hJFPRx3VS4RYZ13oWuhBwUZ4kYMO6MmJ2/g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
A2yt+DBwG6y/gc54ZiwAgseNtZ70OtaReuq8MY68zO6J3zwRWAcEPbNxYY5BdgEGyNqe8sMgYnfo
ZRk2QCy2DIWpyD2voxLrc5HUagO65iCdniOc7uYfBFsYZExVEVF9mXcSxE+MP6/zICOuwe631hJx
GJX4kNwXAblmydmyioWCwaLms/O+ZsNpy38jsrLtp9i1TXovmBEbu1kDZ7dXKc4XNJjABeY0px0G
ZjA+dhtLnSmPWkxQwMpFecckbEHHNkWXDp00gnAciRvK/yZeFRWvRoD7AlKlJXfixHVl8nt5w+sF
0xQ4A5FC8nEihrM3jaW6a0wQWUBmseh69aCDgSfSlfE+rLwf9ZaqbS6+JINp8Soj/9ilordl79fT
sVfShggOfNhQmIIughTstmV3NfOReQQuHLJnk6+1Nk75GnltGV1vTPOTlIUqQgLZxdD8T3tsxVGq
NNeJ7FmHzNiDbLLm28XPgQobBRhF5Df0hihNaHQrKutT2prwoKNHLiOsQIAfFmJzoq6vxso5pCn+
Dg9zmgfkZWX72vkFKDBsvxcGp/lImXCJxLT6xkpg7hM7NepjCma9ce7VMHDwAxBWKMPpftKvrlb6
dlbv1eTf11kXuZm98BSoK8cWwyLvdRW7ntEWT0oG0CKyAq3aH8/2urYKKoNh5ID2VGzLLCcThdH+
3AN+savdnyxHX3T/Lb5KMbCORNzo7um78rRLvAwut/pwA4PZiYOXMTx0ZLDCZr98+CQ0Xa59L4ak
S4XnRXU6qNC3QP6YLVl3HSvRLMxI4PjM8eaPVBI4wI6cYvyTjUafCSMoz5QfJBI2KYuM4OCIQCe7
WjC3mrnLNr1rPQo9ctt7JaPW8/ZZaynFt3lIfbUt8pYyS8PELNRc0o2ikS8sgSPDB6LukQ7deVBu
C5KEQgTIYUwHyKxUrJOIsZnx0N9K0cTmTa2QBYTmXW8GVqwsyRcHosnP6bo0wgIQ8k+w1S1UTkEv
3zhGUL3V2uEMncjsTsMDnyPd8qv/i5Q3PDXWD0v7w/QKlpL3h7ImKw/7uXsgnHbfXAnubedIjn6I
qLYHovfc+jX1wN4fBjHqnvZjxHdnp5mNedlL8mJ9TfT9b79C8vO4mZ7rAt/ok13+EiO6wbBxYkSN
PriQRyikFNlJRRLRsUrD+U1rtvTcGKifcQag0loVGTACXq+d71oE9Ej2uQtNNtGJFKdB0Bwvcj0S
1UklE3MUqwP03dixP2ih0nMrEVaKCLsUAFyn5izJsMIlOvifrcN1bIU239yMMHD0uGrZheIe8o+A
hWr4+W87OUSshP2/UgNIeVFXNfxKbCFnlv1XPxmGuXYHKr4II5T7dMylu49Xs65ekeZ+AbZ/ShxS
3ldcDDO51xXVHY6apZ+YMjOmgT3IAwmkP4yDjG+t3+u0BpheRCBoAPhR5JnwloFJ0otvjdj8WOr7
fU18xLyEPQ8fi893nNQBKYrqBqoBTRiix7f4N/xvTF67xmzxcz9CKeYca9HSIOSbILDoGNBKsXao
vHp+5zNrQ2YYRmIPqKQUFzrL9kt8RCbzqAwZLFNH6kUxlpjNksixPXC0LU4lb4P0ZkGsEbtKVcFX
Igi/Olm48s/SCm+Q0EuDlEm3nSnJjuoF602bXTjdtBWMmbfF2yXjMFtoUeMC7BpuQb0Cj1B/hXkF
US9O17lDbi34OiNBuGqd0QK+DSvJrYnEvE6jZIEkHj/7C8Q8A4H+Cw8jZIbdEQGt1/S+qOu/o0zu
oK6Qr/ECihA6krvj4k6e0Y5QzithdVBFLK7LJH2eeHAga0i4Kk4z3aNh/zVZvvTcpwEfITHNPs5U
+ib0exxYOziO9X63U5b3Xi/F+6laRDVQ2XTc41gEyEzAfZKjPqztV6j8tLnuimZo31TdR1EPwBil
yXI30XlGnOkQCCz4vF81ifIlVgXwo6iovDBqzOzVgOzyUhaYWfAMCyI1QhYdGCqpq6bCvVRQq0We
hnQ7s/WC545Mu/pjcOuO8i8CEyt26vY0bNvplVzUE7+PuGgHw1BGqWBffUXInwKjmotDInhy3qGu
UH998WHIn9jNxNgwg4l+3+k69wL/yxPFyowxujNROlu8xqjJwQ0nq7yT/iP9co/fE1wgY05CpbUi
90yAt3KdQMvBxmey8/uUdBoGl7zx3hlSpvjMSswO3erzrgdwPw1317ZlzS21u6mtrU75o0Uq86jb
tqB90G7xzM6Q92u0iDIf3sRXuxFWGfwdmILF011MSTPR6R2C3lr//B+YQ7BJcYO+22dEhennofBa
uanYql+2GKuxG8hObuZoEF06j15KEuzgF1WG0n8oUzG0XwIaqzp/caS49HBgl7Gje22LV83L58U6
73zr5R8yhoYLVGWv5jQv3q0IZZ6pIQTtOdCNf+Xr83pS8doybki2pKF9/1nPtLzZRi7aCy9fRtkR
TQ66bWrq45nI+IiMYnTd6Mb8iYPjktYyb62NE0uYND/TEVK8EeGGCPhm2xiGM0FE2Qwy2WfOm7QM
5qzjuMDy5CB5qjaYaHW0AMcV1oNQ1vM9usijZKuddHmTOxGfwjoS66UF7ow84kNlFdjaiDOsG863
0YaXZeRAN3yjBx/0QAdEFnpkKBqliE1Us1oudmT8J6QXSL18UA6JPSdmwA4b/A3eqwnWdZt+sVii
5vHeEFiv0sACiqdlPRLwVGGInW6Vo8etw+nI6uY1m4HLscCaZaFv0zuLQKCV8W5c1Ve0dIUMCnOF
POq6Nbt4R2+5qz/ZAYztC0s5vrKC0SF6D3a1LZYeRWFwHXUCD4Eqv2PKiiHoU8VtQD5FPLmy1oy6
K/BL4flQpSA1JUMf81XqE4qPrz7t383X5p3NPntgQ3IcoZ0zG6jakuOb8ocBpf/ARkh7IxCSeNe2
ToGIfIj+iRyQyghz31Go2SD/MWBQ59rAaywf30WXq1LXoaKWE7n9umYwGUIn9EnOLBBn3oWjGeZj
gq2cHr9vkJvPT3hFfBX5e6oWKwqsRv56sWDey3ucydAbwGJTKSVu/OupLK0ziYyRBWfZ3OLGiJaC
a6wpLoZjYs0BhB5Z+FyKahm/yxjYxpwDWxC3kajPe2GPr3m/CCaJTlSLQk/2MQDWVr8siTJ25xfh
FnqI7w+bjz4lWKpaH0MDRMZ4jgiDH/6B+8/PAU2/hRNDIO5Wzl2h06aH/bsGibdF/jLmZiBiQip6
/ikuSarE9pL18J5pry3QN/vJ0s+WBiPTScHJtP+sk9i1aOtst7SrZW/7VPawi/q6CbKxzalW4YrI
xsC2jNyiQx72zQO0nJGDKYGJUGLnQd2oSHBpnGD1f/1xVWIYh+tK1e0efWQlweX1AfZOVKzUahSk
Q8mHuS3egG+OZmYKKCu46C9a/So6hheyYmafP8W+ZJ/7cTxEM6y+I01CpPwwW658+iPkAGb6Ju2w
icRI/XtQnsJrRiWLxR/f9ZHh8WS8cAvYVhXe/plnAc86GPdYW1ov38jA4yk9qozaMmdpdc8IrT+F
ppzWC52xoLUqV6xMb//kxtoTKEsAJYeN34xiQGONMEqppft8jDl2DozCF9eAqBnYmhVjFU6+F4oj
SUA+GUb5eQ8x889fqyKhg9xwZiytAj7llvo8a9BVnHUAqBsrcudlDG+KEVCUxJ6UOBQJiy5/vzxm
vP+FOYFU7JjaCPzBfQJJ0iYWZG08AWDDH3MZi+z/8nf1bsO4AhGOCzmQV+4X3Pa9jJyk9jYZTPVu
GV4Iqxv8SFwIpoATT8i/KaG7Ii7xwUGEFyacR0ngA/F6Jc1aCqFDcifrsM34UVQ+gYABUs7JLV5j
mn4+/uOdzXQX60cnLSohWDsGACdT8WapDTfdszJqIOdkK6QTlWQsy/Vuz0QXQ3prRDgtUTHD38yu
uq8YD2EalC8iygAZbtO8kNJR0KuTEvYGnytW6vgHTFFfbccbkPsChzTvjiW2KYTGV+b4RehLCppu
BuK7AGnXeJp0YqxkBhr7EtRqkcSHq8fTwvexYuCJsa00itNtqsz3vThMOvNo8FLZ/jXHdACUIBV9
Xclk1XbUQVzM9I02oniqzjE96wSI3xY44jCrD1LlLmwArbCktP7+watvhUyhZSqZC4IKBeJAyVFT
GzI/z2hBSvZGKpqxuRCFb1H6vsbTjiMclS9mG4zGQ1y500Um4B3ShcADzl9sHc3f62bFyCVoeEqF
9smk1XZZQMFy5fvh3b5g699F1mu09K/yU8CU545w4n/oADz2pwH+PpJ10NbgTzeGjzvLk68r0o7s
eHyERrpjifh5y5vb//PyWF/gXyMkpjrl5hmkALQDo/exqEPqkz5F+IMtzWAkgkmssG0sRT+Z56WI
akQXa0qeym1gyQ9jd2PODKwqG/VtVSIweR95Cu4cKC6bdaUw2pPGFusjQnYJxDqTzLLaFU5XK9FB
QXNSpAaFQvD5pFhMb1xvEYMDnAOwJJu8CfiqrJaJpWztwCRBdjCrqzjGK47G1D3xVYl5vDAqqdr5
lnbe18nmuNlhozUSva1Gx4Fe/F/TaNFP3BQrWZ1hdizWaKCFzyVK3ezdjGm4yhGwOgZZPEkSCGl5
SeK2O3ds9PXJvu/aU9jO46FEhwVXrxoIRE7nU/Jpw+w51kj1yv5jYBD+eHYJTPb1F+uX6SPOOD5C
twHFFNYgoQJpQ+WbYAZQxErwssXAiMC+g4pUFVtct2tCTHzf/794AqCEtgREx4phoZ1AtIHjW4UX
nLm9q9WtQgSiQtjeo9z6P/tr3KCogeF4J1ld+1csDZC51B5YwtH5aGkKs+BDpK3e7ZKCcWNOrQdo
6lC0y3k4EixjqAzmXtO4EaBSVx/ml5904TrbTK1IzUF9zqtZCSoyK061l5JOvooWBMI3rClJVGKW
YEy2RymTn6TwQqV0F9TZx6/xhcz1BBYDRlwgK6XyRAe3uUsETc8bEqT/YwKQ95KQEUF+Uvf9goN7
qwfMmnYGHGTnvfpDSx6MaqTZ6OC9AreemU4XJaL4UQ9xRmlyzUSMsjR9u7A+6dPVeooEtKr1aHoQ
uAMt1EDhwHch88q0RTukO5fZzQ45rnHNLXlgeFOk5lYTjk5PpQweZ/4R+t7zEW/XI/lwH3fby6eR
IRoK0qoyqQ8j73FpqMM7NLCo5XJD6s4XE/Auq0hJB7SAEGJLO0MpMkV5M2MgdQd6BBGDzXm41jRc
XONe2u24gAqn+O4PSjMBTTYgrqAlxh8vGRipobSARCo4a2UWVLI2JKDpT2Wj5F8ltkeTyo3svzST
RK0EHsNeMsI1u3gpNq5ALRRfLoEH2V8/dRGsVVkoUpnYejjiAWsDA0dLbhgn8q1k08jtIdnHh6dD
VexvQuC96kTcATMC1KegKe9wJ10JmLoWihnhoHY421NB1otzV/iw0sKtVG/B2RKwEBuvDzrRmgBZ
aMKZfaMFHAcVbIQmbVT46kgQ+/mHmfFNVm1GJ9Xm+1WCrlkNru0B6VOaaWZNT/7y8uycOPrteTah
ZrsYM9fGEvxV9zzHmxF/3Nk/gmp1AYwTz8VygceDDZhPBBzHObsT/mfB33GC/jtq2nk91ZiwktW2
DS/N0ItIihS7PEg+zZL8RR2/WiM4TyZ365LQc84McuJOeh98/nXyQcPtmBXrP3MnnA5YxCfQdR/q
PfDrtPNYR/5agC1YlaS4y7wE8LvJB/tTYL9jN3m/8J0LCZjoPS6I+5Gg+xeaAlInt8wmUGoD+a4g
ijX988M8uOlYARO3j9IxaT5opwGLRZ/O7jV/T16zniDEsnQaC390YKrj8eO4e3yWsxjtNJhUkk/n
1+Plw5ScVhwq0Pk0/WSNPhs0ox7daOrCOb3DPzxtaUu6xD3bbS/0YrXc0dz1dcTzT0l/Xf2ZCXp+
cI/rXc3yatVT2dBK2yc6m629eKZNgp0PibwHSgt+qAXds7VeRXqfEiLShLQgC0ZVXVHG+88MhPJ0
lNMG4EGFyJ9E67yRBMlWdmSwB/LUvWSY5WuRBDSiwZhAdb3yCvFjsx/h+wldo9Cr4lrFwwDFSvnY
jyGqS7Alyc6mmSC3F00GmXNGxEeiAablHNclyHdLuvvHtdyPS5D2b00why63yBxJ6Hz+Y/to44rL
QbTj8dAbL3X8IiMG5y8JO7vcQNVaEDg9EaAIK0kmJ2TzpwdKVeXGdeP0JaHdWS6Ux926p3Iuq7i8
vuZw821EoMnSof3nBxMpA4NuC+n2H5/MH2RX4T56cgVePEomZ9f3/udjADNNz47t4ABQaIDZVRfs
vTbsL4iTaYhS6u7rkm9aDXB8v0EO8qclNZTk98R90JiR8b/owYlPNTylOUQkyDzVGtsKF4hSjNtX
ZoiZZF1U9UYFqk6zxms80bNLtL9g6U3t/67cd8USrF6sS0Xz2ot2ji1WekLhUcp1PZJLWHOjL0yc
1yzKmpq9iF38jqC8Cie4MUm+gJe8//TzF5K8z+f3gW3AW6pTX8jraNg3wPWi6eGUZNVeVgF+GR9Y
MC+nWNOvwdOimxizdpY3Gub7UcXC57UeROaKP8L5B8P0YOE899TGOIvFgBNjGouSiRb+iRdtV/pb
YsXu3dsP4AvtopxiRmDi0fG+38+p+FLO7wNz2WIDrmlaHHgfAgYJ6KR1ZilPTjDZJwg2T4n53rJv
9Ec19iF9+sbsxL+4mjrTv21UeeSbPHTqrC9JE0SpXIgn4JOdIYw9uQpF8egHPzwi/8bvO26CXXiq
tAVmZZGm+I3UBuJHy779MZA7T1ErTST9OJu/S7YZYP7Mak35+EoHkxOzgI5besohmgZSLtyvy5K+
yempi7wQOX1/Xg3zEPvgOo56Ukb9JCjo9FyUiXTmYx0VhOiT9LaIgHP+NrAj68SFyngEEiMEWVZz
X0rnlVncXuHDvTr9JOZa9ZQY/va1MDIKjunIWsbWnN+WTY1TwYiwTgp4EHPiP2Nv391w+chLW/Cp
5LIHuRK3oEOkGpVDpbdGdlBg227yTOhUD74VzQx5Yr+mCqcDqf0yXbHtDHTR4FQ+zbv5+IJm5B2T
Sy7J1S/rjwKu/jJs3yUG/+INsVnnBXr7Xo8ev6j9U1SZoZkitAptD/mDzxIpWQaM6f6/tPAO7Q/r
/w+GQp4NzxierFMEd/+Bis6mJC+OCUhYCzgJHi9TmS1rxw2PexG2nxV/icvb0yv/1VrCI1gTilGT
wEkRx6p4ndHhXG4MbuXfHEklNj/q2R4en1OEdJF4WcL7bUtiIpzhwmu6mQNEtD168RLgBVmqHE7R
rpVCV72TAdn3HvFtJZ1dC44UhepMoWNx21+zeCycFgkf6MBx9I1ecRugdkPc7jcLj0msgbq+PqIv
qwKUF7JbfYyzkrk6jpvbC8HX53OG+P+nWOkxQ4wv9KNcg8oQvhLocM4bMhc8+mjNJTCi5H7rRaa0
W6HrE/Bfr7RqY2D4asiLO432zUwGe9E0IjWyVd6y33HyG4WmAB3/xtSbTbujfjFWVZ7lClOuWbpF
ljMLX5oDLyEUNc9dx2A=
`pragma protect end_protected
