// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
MZkTzo9x3sLgIY4Ob8pqU8MB7WbqfbhYGIumziizH19kpRHDEpUFZiBsv/rzFz1O8PP0PhchJu8y
nj++vHU23aSB8au0kky4Gfmp8KEzjFnMP6YJIwPJ63RnXArYhon5hefJJtWNG4ANtX1fwUOhHcG0
Nx15qL1us5hG6J8PHb5O8mTe/j88agVtoi59h7mFvmF//peDIEalIKV7BsF+HS+AwB+jFnnbLoNv
NyZZAo14I6H9DlJ1YDWoNShEQd3cXLjnvQ8oblec/OkWP7u9+iZKLlyuIf+8ud4Px1NJEvI0Juyh
6YGWNAF483k3whsb4yFTHX05ZDPjLvtfA0VYYA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5088)
HjnGcnSrez7ADZ+Jqo/Ww6g10SV8rpft5LLXmyUW6djMrllE3p41OlSMDWgaT1SLvs1/w7rqSosl
DdGGjCZj612e0jkW+nXxidgj1GquNxDtOnKGVNHpSGcElrZKjLoO1LdyKjJHZuPDTpaudeVS2Rfp
2ve5mL90LgMNGHGatXgQbSvkvbA7zsUnX2t0tARxNIF453rpdKSw67M09y+AR/htydL6PzceNQ12
NsCd3cpX1J3lOk9jhaJGA0y9eOU9lTN6/Tv0X2dRuN/bMMo0W6xlqZFiD8d1y255eLlYkUMLjnDa
u/zAXj1L9M0BG+bNffyBBB3YIzf43asuiolmq+maViW2hZ26vOptchxeWsOWko+QWKgRan56K4tg
DdKEaooIhaofJ31b07/yNFmZst394RlwQpQ1p1l7Ln6YMi+W9BrfTurgUWuYmw5tttLZGeZv71u+
JxMJganmSdXnioUi2tN9sgDEB/7YHjz+ipOZfZS7AOPtzDOlHTcYMG2HBXuyDO5iYfwsenYQ440L
D9NLIdI+ZMzVmVL/ytkgJYIBkUFvsbAug5fzq9veaegMmqxAmWMmBcMucM2IRwO8S5hlXaY8GkjQ
Xsk1LzPpNwJWiL8XFVwhwANkXSfMUK2xNNQvV/oeV7Ig1ebYHveAtWe/e7jG5HZ6Ie5acNDIA+8e
wLu+v8qKqatdRSQnGjkzAgA7FwTeXPZRMTGroe5b65e+3/1MeAm3euHZzyIznxr+JXdYGUiZODde
/W2v3dAijUf3p1TR1bziqW1aHsl4C85bL242eW6BAeOeSKKUi6ZVAiPcFtXMOyLyyMDK3ilwMUxz
cj4NXyI7Mt2tc6dqr6XwmqF3hZdQSR7KC82USi53rKi7xZK8Y2S6JhHsg2TtobLuoZwNlUM/OnBs
92qz+rVUfwTs1QUyfkL9GI6OpeEWp+8t+cJusCbCDoFDaXHi44QX11lc8upCP+4egoGmIViSH3JZ
4C/3PY4c2PWPU0z7YCJOR8RqjVby9dcoD7WCG7gwHBnIPWKnZjJV3fonyE/zZhnIBkJ6LQ7WAk1u
Aie0AjwBQXXwl4C6KU6AiNGilcpsRlrzVaiZHIBsu27YikOMIZZ9dyoLoNv7A1W8B8JEAqZ+jxJK
atlF72hJffCGMsmgxiE0H6m37Qs7V+eh5LzWogXtqifE8a4OO9RsbCPIGseK5oii8xZNOhWJRDiB
kNisgj+qY6AjZsNJFQ0CZ8pV9LV8DIWnPB3JYk2PYHNqG4TeIAC6PG+q+56S1k7mk/1rf4EBkA/s
OtT4ieEvHCF+nx7AsJXQQn4q+2iVDu/SDpdsiiw2Z1nA8j41ofzxi/l7BfmK9zxnoUkZOwUi5kAw
GSXoiMNWfplOSV/rcuyk8TQKwKgfh7ImX9WN897+iqHE2qI9y22v4lnjUrKIyGToPcsrPYqKBPq1
GfxXigcrJcKmasc10kXi1egsz1yhg2mXLJG5lUqC1VuS2r8lsCKxhSQD9XSZUqGtzYbFIP/QGK/3
1FvQF6gt2F4qi53IDN5cBFrSZ0CHsYovSTAY7W9WdwNDu63V4Vyh4C5JwDfAkVNdyN9RJxaKIjJv
q/YRTHZUJDq+R5tSVR44+pXwtDckNPw66CFjaTOV93DpqiUkj4S1s/n/kZeMFh7BZajhqY/l8Ar7
btNjAjZ0QhdYYpKCoLFNxLB8+ZRoEPjq2xdzBCZQZKkY2GBPLoWuFWxWXW1t1d0ZsFLld8VI3r2Z
gXteoT5ligY8VkwWYVpKxvLdWaJIov24betQ1dpshjaPFzUx5J66yJSj9u9jXYx8Qkw6I6FwyyWP
+MCkSUc06s0ktuVYozrdRZVNNsplyOnL6nvnNlSw9bcyVp6w6+wOOpTJ4fNAond/hCSgq+rKjszM
Jt1xiYoG8t7leUdBiOIyQe7+SMCq2j24Zh9FruD8FCZepsMGl4dOPHCjfzOX+4E6ngErJ7g0cvQH
NC2dMGTgDG3OS0IC7UPzep9LDoR121fVNiTvNP9o2OF0YUVSkvpLB8w2cXISrJZWstDP6qsxOK0z
MNUEKhZxltF5Zk4HNk6Y78JS3yjpYhBRc84f60KwRaH6xJ2aYG+i76utRlcadsbV5Qv2h856qSqf
A6yv6dtG86wssPnJJRZv43a6Kr1U2ZmTOH2QHfHqAFT0EEoJ4VQvTzq3MSVKPEgEFMUgK0Ruu2O/
l1Ogvy0+CDj/YxTC8dG8l3Lm6HElIbOjWLgy6thQqlWyr2mTNmqicszQaJBO6VOs8kmwPwHMsN0N
2TCaCxA/yskQpAD+WD+cfQ12Rn/F9UQJhpCGnv6QkD2o+aTlHFWxiyTbhooH8SXZlnV5UeAxdHnV
A5COJ/1UWeZhJo5vpFWsK3HWd/q3lG8G2aRqA/KUMcwP4wXEhL1fICk2i+2kEcXGDl0h1L8FXOs1
3cPyWUdrEWIH+UmSicTlY/VPKWPNMqjEherQdWW9Bw8x4RLO0UT1jHJglPIjTvs33lVDb5TGQGCc
hN1DrPmi8pG0ZFAGay7Glm36uLxu1yXIcKxM+aWoQkMzk/dLQkoR/Px3ny8CexJAOw0l3gYgSv7C
Ehk0BX2y7Jpm7ROZJmo6OiSUVdz8hpLHPVWsI4e6GAMPuD6F2w7r+4Sy6RIZz8t3xw3ozqz9tnSo
ZiZM6VR2CHPDZQ1I9XFC2QKNeKg42IQWrg9sOnhTuizu8Vb3fpyEk1XerZRAv1xslNvkTmdKTu1M
TkrJeF1i2BCCiRrEfA7ZZUC3H/UPrXQJuwY5vqYPfZ+Ra1YFeYwO43lkfgtOZsuPw1jFZJSHb0qN
GNMlxDvV1UVmDmnNi4uVDKOhn/fsOyjnntAAvj0bXDQTlqkzII6HUQXn+LxZkDJVV25jJoY0F6m5
DJ8n96aezE17vbt3tUkOGFJgp4UpuT3sWd2iXlsEfaUEezC8lFVAluFvudgJWVDkICCU8kMmwgHi
f31s7xyByfp4vSKhkOVaW9aWjFC4kUV5hPf3aTzEkUAbtnBDhF3g+AG8DoKZwiL4UDEhKr2qiIga
kdKhcse2VmtmRlxlUZF7sUnFKBjYjZeeSYanFVFMdF3SiJg4+rr2dA7hUCfiI9qN3ZVuMtos/Rrs
wT/c8Ea87fsnARPlHHVWQu3SbEXKn5pnbK6sfQEZaUtT8JvY5zZNp7OMpO6Exd9N7Jnfz+iaw9Yf
UTd7NoC/n7VruzF1bjTgl/mfJC9I2uQNmGoQnPvNOcRXkqKSg0jjJLRSoPKY5OB86aDGda8zxBSh
u2truCCVxpYmEbUKJr7CDumKiI6wlk1K4JgAM+tmPSqa3nMxgmzqF/xGR9gGekIT4PVVXHswlzC2
zcqpj0fEj77vK2qqfZb7rWe3Ro4hOhroywGIlYCilB4AI/KXvbOajH2TJ66FDbsU50o7kzINHZFn
ahSe5Ta87xT5RoGn0k+Enh7untFwWnu397aqlzbKy1Odza8kLqt2DAFc54gZk9Xpe8K2YME8yn6h
ihxS6nemX/5+UEQn1zM6Kk5zbgsZYv7mxkTWhl6WlX/Jtgr02Y2C8AzwKAp/lcys1RqGNGZLuWIk
vaoZq3mbEWeRDCzbRrF1Usi9KYCvUd6RThiwnyG8rBZMd/8dAUuiGJCE2jiDM0Q9syy3V0CHM9i1
SCzVbs5xWGkj+NioX3PgaxkUzCn2CBGruhl5xMhmz1G630X9LDlkqImMvh81qwnf/TO7yTgRkvXe
je+0Qa6hGbDMy32MD8d4jKsoWADcNs1RS5pQ3tkUEzm3z1bUYhPMZtSf25wrlVSJgUHnyaDBu+GT
Y4j9eZ9x2eZfEPCUM/D/6ObchvcM8MWyZtlWQPEBqfNOnUb7fe+iaFDufId1Ik1y5kgC32Z/+oBM
b8mZXq7XBac62PU9jTqwFfn6S/Z/g687gLemiPPFU8OcG7E1PnzypsgOeIgaWFYVrQ0lh1zWodB6
DQKltyLVc/iC1myxx5ZIO451VejmWnUhZt+VCXrGIf4D6jPY1oyzGkyfy7mHQ5gcDOeTK35nTC+a
D6PTob/m7A5MYZUzI3NAOVLKG9vDvg05NKWL1FYgoalBZGpSCZI8quVE7f+RXC7y0NV6E5WZak8P
aef4mdN11CLTT94EqIe9iFdZM5c8LF5t7JebKImlapRz/QQU/+cp7ek40MvMRveSuwgw+qStdhtI
q/hSZ6faBG559wiLPuZy3Q0jM6naPmo6Zk9JkjpRKtvRiP+X+se9ilGpLhSXYk2gbuIU88ly4TGd
CYdxCowYgNonXo0mSw/ZMDZagYAxDG4lpGo0b2eFoLm5BsPgJlZOpjtWgjvGOmrQmQAeI9lzUu/X
hOL9D2GEI4OuQoIcHy8gjkx/V1cf9hZxQULbxfSSxLUcc8qsr98ilYZ4M4jjgTzXz/NMvAgDkAM2
V6nN9zp7nU+D3ayA/nWEwUuvF1AqBzQKE9DuFxtOHtt9sdKEIt1/4bcxmFb0552eFp0h//akl8ns
+4V3joBCl4ne5EONZ633DWzUg4NzoTOodMIoFw/us0YMfx1pIRO5mmnn3HkwyKDnWsZsUVJKfLtM
PBItKHNgGyHnkOuc0gdOqSxdJy+5e6eU1OJG71AIT9yQ3RbOaAD1wVV/Y2/eYDC/tz7W7Dk4pBxn
JKjACmycAD+DxaTrcHsjTBLvNETH4o8+O5rV7lBdPqZueOWe1ZJKeZ0heWe0Q16y6xzKzucWcFf8
364yPUtNujikwSzM9d+HayCu0XH2PyNbCCQeBPuwv5K449VvSXDySPWIYg/1W0cd7+Awau3vJZZk
x8j5YVnZb3yiySdgkKGyKNfv5+bnaVA1DbI6cnkZxzpAVVvgA+DG5EAEb/r4ngERZ+FPeGOXjbzy
Q2eXrZG3jXfUa9XFPdGB86Y+ac3h8TBIc9N4wxwhjYVVzzHScoIDEyTCoZjIeTDGf3xXZm8pSVG1
rxMDJjKJnAnin3iJT4Tx5wgPn8hDFfgJgCjjfIvstadKkly0hQ5+3K1kcaMWCTFOZtS/TO6TrKql
8+NTSHbCrgWWl3HrJHEy5YAQWp3MRlSNEKwoY6ouOmG1+/54IA4IhY+CriLLZZEY1mENpCR5hhut
DqNMDIUsI9N7c0vWPO2NOlmbEdeY7ZBCSIlHFVkh48ZL2EnSclVuaKH2v7u/Zvk40lgOwK0kU4hD
bErbXz9271/YyANu0DxKSFs1mu43N0h1I5hN3intESUaEUPmaG3bYBiYHGpGTOlYS27BjwLn2gkv
nGc/EfAZpTeZPq39BWLad8Q9e+M+vEQP3bjUs0xr0k/NjIp3A0t4pfLUWJBGhVj5Bh9LCLMQXdCf
cixI0+FHTn0aDtGIxyW9LA0dYY7dYws5IdPE15iBHIccJ+ZF6/ozq6BlToMHdtGdYwhiJBVJVo37
pHkmLg0vWlyvOUSOB+vudRKKTHwBBtzb8UUxEQ3nmVS8N4ZFRe3YQvxtNOczOtUqfipwlixc23yY
RvbKYtWu1ugFq4tN/uUjxo7oWJcUevQck4Gu3L92N6uclFxJVZWmIs1RIvTzOx0Ymn3+4Yq9zGnc
LHdcF7HAAEDoagQ5MAXINuQ2ytBbLpgG3R6iB+9IVxcUQJnVH942kgXdnG3UCT+6Yx9nG/bOhKp7
+STG1AYxxrbAvBAVFajXtbGMdOPstvXyg0mcVQ4ZsbhMZpO46n+kaN1RV7KQenjbOQu6/H9W7DYI
DB0UJeWmy5LRXUf9aWiiLXyUzAcP3dGBS4o7gwh8EfwBlIUZXrhUq9MruvuuJAfQ72f5iaOZMla3
Pe/9MQK7JkLpGjJ9phapEKBzbN/0eS96PluUmXYruWDaiDGi0Ict94FXXB+WoJ0hVLRz6x81KISL
9CEVWMFDuKTIOr00/HdoryuzEO7UquAwAzB3YoUEP4XL+AqKK9lcbW4rg25/fk7Iq5QAczpyvLVa
5nJ2PAHOJAV1EqIJgAcrFGLRZ2v1csHsklQ8uICrm6TAcNG9GbhuS8nnZ8suh/tNvikf96DEsrJ4
osTU56P6JdCLd+ZzOf9qavIsP8/XvvFMKeEWVFM2G517ItVq9yMm/5tQccSv9NZ132AmTJO1e2CT
k2qWuCFrfe/wWtK78JfMydP4bmU+r+nh6f9Ax/FNs+ITDrOs+ZsdrlXlvitugV1QJ+Y009jb9iux
kFO4dtV2jIXqOESfmfPSNO7YV5GTbeM+GBmPPwIHLP3nJJ2knpdxB7VVYfYVQh/GVgIdgy4gM4AX
zkphxNCt8HzMbBW8TJM4McCgIRpLHuRwMoa7KtgYh4sk0QIGbBDNQmodY9DtLOc3TlGItR77w98Z
Yuj9kxrzbIAcgax1p+roUU60RLLQ50SxFADaOuWBrLlCJ+trxhbhb0ZPsux9exRI/VLL3qaN2cS2
sGS+hWtBEzjIpiY6Ycarpkk3OPNiQB3DuNwu2bxrAUwMz2XtZLqz2azoxPFonOF09WukWqt7oNB7
BHVbZJWsg00xayiOoXXJTUwi2mPuAy2q8qq0WS/osw89/Lppaou7lnC3Nn/t5plzd31M5X2jbiy+
xJaUltgOgJYTKNGyUzWIW3/bKBctjilnGYJorMFDQSdg2Kh9ESEjSqUW6HqSQ8kjvhJ7j8AVF3pW
+TiIhpC5KxqO/HSn+IzAtXKW9ogQEKad3rIaLjSrl0xhWtLPwftJod+j5JaipemHwYswOWfUlV4u
AXNFDEGzedB8Htj7+sk2jOrK32yfGnKG2aWmSY4YfL1Z/d/TLNL2lDXyvIZpTG/eJuQgTEVicO1k
E6vR2broUtCVzer2DnfB
`pragma protect end_protected
