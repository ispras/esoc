// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
hFKupALrMttFmtvG+wWFQnrN99ptFTsfUcwE3yOm8t/qYEibAoxbag0MvqIeFPlV
E2LQ/oyG2biJ6X4jdzGMulvyxKB+lwqZ9K67G8WVc3YnyYzmu8DQPdRTTYvtfFAo
DDyZz0A9n2tnCDqhZ7qUrqAhsrOMIvKK2JI/kXi+y0Kgs6KitF7Agw==
//pragma protect end_key_block
//pragma protect digest_block
SIBcm8sDlJOeSxI9TyacNjp7Qj8=
//pragma protect end_digest_block
//pragma protect data_block
hca0EhxQi/EkZmQhXI8xGQs6iB4fK8hfI+pKDac74Zzo/Xg9SsxFV7nYGZ9PWh6j
w5qSiQt+qYBTXgevpOKEJ72rpEDAgfR1D5CLC2MYZmnT0rORTHfv25uAM/zoECrX
R4kHgwX4f0s+QuLUfs4kr/gH3GRvM4qijOtdQiiyrSaEY3bew+kqu2w/shJ0mW6i
wQxFTJvw2lTiL4RwuHu9KZi9pnuwF7WWIoEPhn5W1ej6Ai8rMHF6c/0jDqETkYAx
MOkn9RLo0gW6IDbKa79NotfhSH9Gx40VTM7HV/DBCFpd71uZqUsRH0KmK5jd/5o3
Ktz9bEXs3GHP/g0w4+cTdtBb2gRERqPWhYeL3wjkERP+C0GazkiVbnDx1GAE57hy
lD+IRIlVAABIpKBsEkDWZK123xzIsMl5W1gusBBoNeMDbrjuP0vD0erdkn284IXm
WXHSIYhaCcTQNIlEyqUgdekF+ODJtzFrPjsaP1wYvDEwbxuKMb9WZIud8zHPbgR6
MOquq3etnYrSxjYxNqmyPhb/RbLQ1dMRjjt4FaPByLQBUn23qxLoRllQoDZC02j2
SSc6nSa6z9BeScc9qgBYocn1wcEKoS+kkeOsBSkooq+9LfgYuXHtTP+NOx5EIEJK
wisB3H/urgEUttvzSDx7Xo8VrNKwxD7S7+eR2EUY0+Oo48Um2ttBiLY593lzom0v
1iFfqKI8PhLOj+eBgOiB5ytSsBPDWU+udrzv092+RDJmsXicqsCf9IHvFofOwmxU
Hw+xeISqJi27ICPcvgcLs3pJHKmyub74KFarPKlpkDy3t5gVlFmdsW1BAvqCaWXa
gVgGmQn7LKKT5UKx//mSkEiW/KGfmOhRd9Dz4H9ksVxsM/ZEPpiaTGMiab+nOiaE
W9IiGfcoNdofgwKP2b31jnuWAC/KFv3guVG2sW662OkZn/C6JTExk5hGNLpEaBdy
oeyfSKD3X6+boOB1D5aZCASvI1GfPcGVdeWXW07VRcBIrLGDF9Y77X/YQNJPNQok
2X7Ky9SSLy/XyPNdv95jpPo+OqAefFljIXeYkzWMeStQmErKe4g9Bbz3vgWvOS3X
WrYismiO1Jwcmo7PAqs4Lh9nfcQqu4UwrBPcDjX1ybzh5R6DBeWbYWZQC6J/4AsM
1mQsOxEYPDFd5yXsxcqUHFYO6dwka/YCWKQkiC3bM6RE8VSP1x8GWhHopvCM8tu8
C0upn3WaG1mHrxjEcFclrnycelt3Ceq/jJb/2eZF/2qSjqczg3SqBfxRAhmuVkiL
0Kp+a5gEnLp23G5g7GyBIavSS+qW0LxouDn9rjugKXDAJ1YNkeMoZVJs3A/sIuP9
qyE9l1GuZjuKhQq9kuvF0pnL3HGUfKr83HJfepiYFQBOI6F8N2ZajB3VCUgYFSVp
63SnAKwKP4IuX1pKJSCa17OCO1tBZ28sTa+Fb6wewdGMzwhtPB+tqGXSYh/mPCEl
2whGwUXbKv/+serIrMLyG6/aNi6HbufaRfUbqtH+Lw0eyd1MV4sGIUAZM0NtA0Fa
KbbN+bXqvAJmKV/RzrfuFzyYLMzRodhwIBc6hLD9P7uk6hj/+lrTfl3nHNZnprFa
wUMDtxKy54HywMCXneYdcnKtsSP1sqNSku/Ouu8wZGkEuyF8pEC3DrO+cVqFmPKe
yu7agMX9o9IqZl4aTz2llKYQRY+r5TGAfPdIhfpBGce0WhhemUHBKQYm7741S8vu
rRkL29AkRTQOaTCHIgakA/Hbpc+K2NyYANojjltCME1y8Gj2kW7ee3/+tf/J1kZf
XFMxjvjO4ljgRPThWs/rrGFxfUFYlIG4H+j7yay/jLAFNfEj8mSr1ikqrYw9Yqpi
OCX8bnGEdS1pd0bHQW3EF0D5XYI7H2Qy6KyZD+/MEyoB+u1+pzDPqGIusVcq1Tp5
wrtIEVMW2pwgyLsztq9BXhbEZjvthNmn2NsjuCAWqoM2OV3Y9d2W5dp6WrBoinkF
nS+aIq35pjVOeh/dWjz18yIzyU5Is5xwYGhwdDmJbx5Pn5l0X/SeDXaTsTYvORs0
lXZ+gzwEBMRbTWV6rGhvjQYVspmXRUjgwgHNpR+lHZi4a8DZAutCLWZMJgu0kkhR
boMBBLkgqNf1+5GxM12bhnmhRQIqOkjNZYQU0ps4kXukX1hikHVsoswhPO5GSxv8
Y1MDWmYPt/VK2CrjCJzBtyQMciWQ3dbj9NKeIWNNVr7o9I6rR4zm0VPlWr2PznE0
nHUm9s0roQ+6NRnuyjziX3srfqpxEMDJKNc0qpcf9YEImfisUs6Ha0aGfuX/gyHH
N/5URbtpSpuiEEhdwWs5SC7j9p1yGpDYevuZ9kepFB9q8Olhs6aEf/aqjkRFos3y
6Mg7QDg2Smh7k37pF9OIyAjltHZa3HK2KJWa/UNG6aF6sb8BL+uaGqDvgkmlGPbS
MB62tr3rw6jEUS3WgCCbIMPhheChhIKGm16BUgbtBwtVm2AOhDVBN7k06oUAcEMV
6Xx6CUMAYrfzUN0SOLQzrDgFPfNDXy1SU2U+8GoYKu5lrjbyiOxVcbAeEC4HNhTW
JZ+hQu/lc/SFBATCNu7MnGn1ZPSUV6/OMQez+2J+ws+5QNAk77Q4kg3IVM9spLtL
0Ei+g4ObDNnitRfVYMwSVJk9ksdpGB+WV+Axxc7yHmaUA2pdJDmJTmuBnSbzcO1z
VaYQe/kBaL81lmUqhiWzDLE3WQuLUdVFTa0nzsc4ATN+kc1IfFmEQE3g3Ld8oRst
ZIIi8cOCbWvNubXaKgIyKlHUxiD3g/dHvh3KCkOAaamwod9pxaOS6AijRHQxLAbP
exDb0wRG8pfjyFJYI344wru+aW4uAn9dFe++huTw27uoVO/3Fh3MmitG18iDpfej
sKzPn3HP3OCZ7zMc6Gh6FcjyoLT3bvi4G6xh1DdyaJ0l3dN6JM1BNopzMI/R4+gj
PYgk8cU7vYXe99GWaonqVpEJbp0+6ocf77F3Qjo3gayAQ9V/QHOj0V9pCGIRumnW
jIup6Sd9OQcGGu0KmrFKHlnTu+tc8lJ3CzQjkOcndsjV2yx88KPqv4QcHlwUItWh
tG0ROmKU58JJHRNjXq6KC0wmqU34kngxozD/QvLRyDmNUdFHvCvM9AwBm0wIyvNm
34oQ4OabRN4/CUY92VimvyMQsclOXoU0TosDtBxY7YuUWEJcWmRlmn7Z4shc3/aX
3+ougT6ziJVUu+Gzwbh/s+gdL+YwMgbelxquEjn3YoSmaJyVcubBw+R3TAMQiFr9
fLMciHIJG/1MCBI6M2EuvnSyBdKmCZaVLT0dRv38gftvPHnp6elZa8Z2aEAk8DJw
BJtOrMVmK6/5pYn3moOdJlg/edo/Lqlh9cTDkW1Mpf7ejWKPsMlHnJDL/PPDuovi
PWXn2MtgJbkc7h5LgWnKE3AFKfhXpmS2ODjNL8BZnF5QkKRa8sSSxXQ66H+ocjsO
1NSWmbm4smQK4WwnQDgY2r5L2XfZjYb6Mdj0UjRRa42nRnei+tgxYv/w90ebSLi/
vXTwJ5mXhqT/heAizzSvPy3SqhWfXirDmL0dRH3KXV7v9bWI/W+WpTj5bJxmJuuC
Sf9VrPMrx3GJHyXFe3QHIWvMxLYxceQ8SOMrxLrFWjnYVH+kukB5VD1WVI5y4i/7
DWqp5zJy/I1vDbZE1tHBpBNDMkAG8TAPJ18IXvH4EiXAOmIS48yYkDLKjTGUe0ki
oGyFkHfYNdIQ9Kk2bxDOQa2nGRxw41BHdeDJ2XucYraqX+WfAeaN6ZkLpkJofO/P
Jdr0H4hyRlc+bfZ+IokVnHAc/osKUKIiDdCt058+83RQUeBIPpHpIgOcmVrfvfsK
2vc2jXd9P3aUt1+G+UphB1IQ1qV6LSO/KfFEKxawL4Q9KMJobqj1KKoEx2YqsiIY
8Qk78LYsSEe2f7F92dp38MLl1DTxD5mZ1VZOEKT+TAiTBt3wEwbWER1w7gCVzip8
kphQrSyUOhSpvrZtsu194bix4vLcdNfVn9/Eq14I4iWY6Pt/Jl+HnFNdCV39Ahsw
fkVlOTTCDPPqWCY7509jqdjo9N+UCV04ezXvkprH3cPuuvV9pTdi3MFNqpTc/tx7
4HxtcSnpMV0wXmzuv1HNLZSx6A4havH9tUrrrf1ZE7BczWtHYUhknKqSFM2nkF0f
5Jc3qX4dA16RtYzWoVYG4ji+hjreUaeR2+9P/79UbZieHf7ipOl4rSzyLE3r6vvs
qJyPG57WkyFHZ7JhMFKo+yScrfJJE8ZOlmi4BgE7alQVLEkHHpC3tcT+LFJ1SV9o
O4IV0TT8mOaZdNYpbqWaT3XmxnL86eHcd+QhEV5SplEzkwk4TeJLXqoVsfQDdijQ
ubo3Po5Xz0xIHcXeUXOd2IkTTyjnyZVg0ZZSmTmXCFn10EbZh8h215zm0QleWl3t
eNnoSVTLq6k9RPP5yCJLW6NWUNH+9RbXs+PLlH4BeXHEkJVMmeewIuqSB89rEB/4
iH0W3Db6d5pt+YiMeS0r5DAGYOKTwumfstAlEJ86jJ3qV+002cwXcpgr/CucV8Vp
9F2Mlc6CNcGAr7QZfXBYi/1TqHTjcfqhbvBaQMGNuE909yDO61SH7mfub+S7yUca
8nZySbc6vUuzbFExz8xC9Gb3Z2sr5RybIbJ9Askr4k068Ha7ne6iOHiNBlhGiMHJ
pTr8dJxL24OlmGy6ada1OawJvGYXSGklRzpxszm5Kw0osHGMU11YvdSgRkEEtJk9
XMnSCOso9I8h4fqpLZQHRhZL54NaR9/r3OvROvn4JW91Vj5RHoVZjEw8Z6yP3kPc
q7soDuxB+H83Hm/OYcOA2OYr9JMAmXqap39FhJDj3uVsGpn/W8XQ7/uFazA3/RYx
Ce782oK54D2WuKkUDbYkjapxeMRoMMjFXEzMQqhYTaYM3QP5u2Dgyp0obQZRN38N
Fmo/9attuzHjWMkai+HEedEBHhu6Fq3uivdyji/7uVyyZFfxWw5looCGsEb2BzPH
NjWO/vS+YCqjD08HLBKlF708LHJz15lr3A4c2BjW3RLHCWXhuZRp8eCRopNqLWt+
u1MIrulHzOw5nKKR6qcxa10bdYOBi5ukwxkuRuehwX2cAuJnOW0mT6aVsijR4O/E
FyP9oN0cu/SGSOBYC965+pXF+nICQBPl9Yr25iXPG76kRPOntxP9YgsQ3oKcHr/R
Hr2fJvIOCLjAPZ1czwXLbjXT+VDFdSLVw3jhfR5qmIVvG9VviOfPW48uCsX3teSC
VIXUY9UG8mWtenm3FF/4nXDelw1zouVeJl73d2jh+RfAgt6/LsusuWkgJZQyaKMU
wX1AGY+GOKpW5luyXYeDIGoyF9Xh+FwrxqSHveXZ26hT+dOJa4sh8I0DSgSY8Pc2
lBzSU0jRCJGt38omjS8jaLAtlaiPADg1bkKzLa6vDh6TObc4E8m0HIRLERXiHusa
DXUH+MK/6DVYt0NcJsSkpxZFMF7QvuRJtvraZsU3yE+GJEREz1fMPTQFleoJCnJa
Rdm6mq5cLqoZdxWgv8/YXz4zkDydGwbVAmGFuVcXDygOV/5BEuInEtns+xqfeiE8
axHQ6x2FKAezuWhDlarrG/472+oWMAKdbWu8ADTHwwt8fgHnsAtt3y3Th/1BhuKB
oU4JsD8HzOidvJeMLeeamk9k2TmNm28k2xp2PDelGRYnBAuYnVs5eEQVUV0CsUgE
2+c6OK1H32CSVe6sksnrUqQdRvD3xipaHHT7EK7/tsSV8UbQO171qK5cE4OCQBAZ
P+DM+M8PzmWOw1QWXhOdxJ91cDq5vO+ALTyeFjynb+LzSapMyTDeujdR1wBP/yzF
Ggmo6J24exiLVq6Jb7ZF5v1DpgpCENSK1+WiRcPWqTK5UkfRYindplW+ZJCCKruL
JkAXsSpfAtyW3n2P8setcFrNFsiQrZh8heZQyYV/T4QBVkMGsyCP8mYoPW5PeRfV
yMyj6gcyp97UJhwNUAHG1dqjnSfAoiN/2xTN7DeLaydf7Fa/Ayzbup52i7cntUtB
yBgzg4dMPK4HhvamFwlkNjWQwet3W7gH+0FbtCt+yhpR1duOzUc/sZHlodHyCdma
fipDXgChkvd/Y3N1xQhd4zMp8CwiBRXWmUTUh7tlp7ParRLJZktqgkBCcEuTNmJb
HI5GOQ0lZWkGKYDWebNVhZ5PUGXy0iqMO7rrQrLZBAe9UgKn1gUHtRxpg03Z2T1P
yEP/p6D+A71JaLySTK2mQW62wWGdNIWj/m+N2VtZe0SVyEnI8QaVrZxHsAF81P9x
MEAJCfzG0V2wzFLiwEA0Qta3ttbzUjOycM/yirKcse5NBCd+I5nqLf/nlOwImQSy
adOOfGkTBc8gcDy3ikpFVMRr0Yty66c7t1xyhgM6SUfTI7RcOzVk5BAOiGr7FHVj
SKBdiQ+Xiu9Ssk2WHLUE9F53lbdTp9WbCP3L7ulV9tbue8mQott5U22MkKmFcqdI
3eBwY320LQmFTiwmu2NdtfRG82xr2kb2RxuAFPzmdh9lKLde3pQN3EHgmDpc2rIB
T+v5FPKksVb9K5JiTya53WvBqstXKKPxHnJ1txNhetQv4ifLp1k0rgLE0Tl/SWTq
x4TG7TnuFLqWg/O37xeLMncAXoeUB4CdMabI0oEVLiiAcUaYk3iefB24RFhJiT+5
2VSWNs+KcWasKrov/X+m5yDxgOuKmDSTJ88aQI9cBKAbkHoun8gog8IFkNSCl9U1
yXteGF/Q4uKeFyIIgFbgYEqOeC+rEWZqK5VBz0RZ5CKm3dUMPZQTe81Tc/XwbN0Y
RtNWAp2NGT0L1jXW0M15TFZV1kCtiGIm2f+Czh1Wc8riO1+wM676bJ0qXqxtxjqJ
L0lUv4K291/LqBvRGOGGmGEbw5ndcnW+Gw9fT9+bfv2BqKsLEHj4h/NR7vT4G3O1
oo2Y8a4klS3tTwWd/s9CYpRQXEuUuoRys63FdFqJzbXV5QG+x1cJ106mypSiW4y4
ZmTSYnPcE8SOOCNDF/v3Y+PQN4mPbDjwDRDA83lcPYmNuyQx+2T4d/35+1lvkmlu
c8VtFy+LOXr+21ZkJa2Z2azo76wEZrTrdooO8lnCfUuJRSOCIP4wOcYB6UTX2Euy
p8HdtlFE8tycEUCbrD1FP9gWmZL4x2hvB6FypsEYFeiTc4+YPew5gohU3CvP/eFZ
taXst53zVNj5OKSBHQ1TlCI68hu5Ba9pvks614BW0KiQyY4rWJsFBveeFTVpm2LC
3Hyv1xeYxfNfJiWE+XvIQsHV71mNY/lzU0Yec8syELOVQTVMpvm35EjsOwvPRF6o
bYwCUVhlITk2X/Timwzgp8tVQoOFNd229P2fuYUVPajxCBnw5LDcbTo/e+bvgcoA
y6clj8/L7W0eNV6PLyYLyjLGGtT2LYfOol67Cps4QzHycXDxDF5/IKtr1YpHWVGg
wLaC+YEvkNdf0tWv4EmYZaUYQGhGKgkouXzOY1CzhtLh6E+jsnd4jdwjQKNx2/b/
hsM/X/xQzpdBH907huTcYiz7WCAVIbEdSl6BFctzgUg+KFKDS42IBlTXsDPBU3DA
9qfmfR3EFyqfkWtkrnLEKX4uaQg9tQFHYGdHsQKUTmATPlpyHx8vqtkmSQi+WqTL
F9O4VhZnFOflZapfZ6QE/sHp7qXDy6m+Xspp/qop96C/zK1TEH5CtEk+Ar0gaxrS
+cY1VN0BL1LiFeUKSjBbxfNCrpz6NVm4jKLe+F8rhsMY0KA5VMNW91fAUnAFN0fU
iZKYTmdTHV2stvvtHwrhnQ==
//pragma protect end_data_block
//pragma protect digest_block
iX/wlKI9gxmE4weCAjNecorF3RY=
//pragma protect end_digest_block
//pragma protect end_protected
