// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WHz81zN9sUlP/8/sWQx9VmIUdwNl1/zMdCF/qbEyPZ+WirXxydWh5XaB+eQFIsOS
RGyFTuY8NmRpEsM2cuyNj2uj+m3AkM2/kz5HehNpNVzTU/SndOZb19crUmM0CG3M
g6HIJUR+3smieGR2GG8pq0T5uBPap/7rlMnlcELCbw0Bc+rJ5KHmqw==
//pragma protect end_key_block
//pragma protect digest_block
G7s/Ei4icBccuYPoVeeCp8ylRUw=
//pragma protect end_digest_block
//pragma protect data_block
Dzf6KZgE/oh96WA74gRdC+DVfzA9NzV20ONls0I6wZYLvCiHyuGkFna9PUmjaBHH
R6noq7LvFWzCRGvc8Myw/Ae4XNN7yLbj0JpLwqWLo5ceUKS8KZQ+J5aqo8oCRTqa
Z8AqpNOr7exlYeFPsk3tm6IFG7B1hWxa2z+/w0iMh6ePbpIkPT3XrfKdj6+Nioxy
uTDIP0+UG+dtOiIbtrB228GvjXC5VPQZk0NYd4jHETfVyO/zR39dzc1kgaXEcbA1
48k2kUY9uzicMpaKcHE12ARcOkxqiMOw6fB8750+6y7E2GBgwwLhbRDUx1Y8Hw/X
Uzjw9de9pTUC0mo+9kPJ/rBSJVzNduk8vsGiP0r+mOsE1fy5yscKCzPxTa/tfWk4
xLypMLf9dgLsg/u4Cl/hIXTJla1hebTHSN1e/WU8I9VgsfuXG+PLZH+P284jH9zA
+/krPkW1g2DpyVLhx65MEH2Es6USeSMMiibMHeQAAw3eQzmjJxX06Ic5XRLB3OYK
yZRKH02+o3xXbmDG8QScMCI9BpEfV9IK3B0tCxKZemvLHutfiC27Aeqz6axnAVlb
eYOLSAo+IKurfYXwmy9s7xlUIQPPTPWqIuifSrvp8M1VqLdMB03oH3qtB5zuBoEH
h5Xea/XaIaDjK+vhJTPo9bVMbQFP3fp3O//pqErmgINag/xIfdQ1VOrh7ITs+avH
n7TRLhLYiYeYSxQnwKEgOMgZ5givw2iz4gFlN7/Od1hW7OHh8Uu5JQkHs2xLBVlg
Z7orJxBcaYbo8K57dMwR5pz/4Xs2MlGA5oE9wnhaO55gK6+XHK/i3oyyXNek5RVZ
DiY43ErM/PvMTUwUkORwBcpjE+cnqritxp7g+G5gd1rfLEsc5/qxbHQ2xt0LaqSr
VKzfM3+xcWVyL8KsWUPibMsM8L/VUitmcgm9xhK+bOLuk21VRydstNoXW4GRPKKB
+IfUwYho2nm1I61FLKh11+iIoo9l/CjrBx02hyHTuMTkIyzNP3yMxpNzD2aRTMk/
YEywgoDfHinBxnhTJPKSAWb1YSBFmpWtZFpehMZL+7By2CLjzQCxbxDqgXQ48O2b
OBKm6Blg+3UOve/nyNOqR1mIaT4qUEfPgN3Sikbz30yBt8ha/llTQ6LqnT0v9yPs
+H0Y/Yr8GkFLARN+uIvhE+GHBa+JjsMm7SKP0j2iGr8JclpQyxTCyX8vq8Fdkq6e
m8K11pVatXUWLY9AYzUAdWlrWguHTkn5+F/TKFMxjw1OtYLraHOv6G81EDv204S4
tPjHKDM0ZIE97Ht43JKlcEgi/RMQdnEoz/cx6CDMdY5IKc9wiN6qHyoH3lccVsYy
1mndtvAtyPlEVM0Oz7vcVP5R+qTuAV1zGxEaDTqrDHSH1QeEeFFRRJk11K5eFu+s
XGwxxJzNwsM0MxDUzvH0jggSjibBn3ciVWAlxWUQzqGSg3ElHH0sTSHwYw7YEXnU
10wPWK9DMzyKvrFH+KnjxBIObJoZRFL6JQEZevfPFGM6rvxc9nZJCwlTCUg120FZ
n3Fjt87di3TJBVd5cKxhRpr/qCUwH82fWEP7CEKox2QTaZC7Pu9ldyCnbQUTMYlP
sLH4oa96lm6pMHkSbVN/MDmokctTHYAZDfEZL1tavRFKtPbT3u79BJxZsTEYH9Jn
T3ggM5xHTf86EDObLWFNdU+e2DuIni51lQqGGXNI7SOD/jp5S+0Yekfe4dz9yWqO
RHZlhM//L4yb4o35hXTF7PjujXuntdd9Mxhj45TFXmLxm25n0aLjZlv0PxbL+q/9
qXoTz2wLl1g2L+yzOjIMLPcrVQ3OT+cDq+70Uw0yjrxDBH4bTVyqGdpOrnPeJc9I
soBhaaklk53M6UPd4TxjR+KeDP4wuK5UyFNyCT7zqwahZbhHEHVKpvelMNXl5vaD
/07iEw9toEbRlgXLRtHfr5/gXLbZ+dN6K6LCDRxsCnx7QziTleK96eHVX4dPFhU3
xacWXhoHjTAXMe+g1JjLpox7elnhJXwtr/CL3p/mxdjBaD5ooo2mn6hsMX1fwvCR
5qDuYz6E5GD0zYDGR93/DRlGfBeXednIfXaVshJTNwLsllNRtDW7W9q6l2a7LxSU
uNoIUwmmQyOfwZ3MtjEYmetMJ1U/DFtkgf+mFgn3fgZOAuMK813BvDxrPx6EVkuL
eAsYUcYrH4cxGlYoe3aV2WruiJtncygDKOhk0uUMdfzgDwT462u+P9lTR6F/8Dcx
gs3gfG3FhaAjfYu1LyPcocw1MpIdFRnJ5U+mvKs2vkcPirQ7uTtvO7os92e4qHEd
y0dBf1hIv3LWaNo12IHtwgZ5zBKwSFkFX0U9LCkpGA7Oey/z76P7hQlJxSwqE9Pd
CjyeKVxCwsJCli7xz/DQo4db2SyPbOwZY2wcddDzJkSSATQGOZk25k84+YfIycK0
AU6QZ2u3RSxqt1RpkRLiPTgynpR57th2rLxRAwCb/oIj87tblXHPVKTD6l6AQg68
bhOnb6JWuP0/dNujWuSGD8eOexvA8PyAQ3o5fN7eRD4z6yrbwmWY4CyMxCZPTEnX
4pmEzjiLejRF7886VEQpI1sguKKM0Gj3+Q2EAiUFjATqlBJjGq2sX16HXzi6V4x6
g658IncVOnb+blsPiTS89Kz3xwkVd15nXbdQ3he9IuAw8KnUk8B3fcFkZaOfZ6+B
SLn/IUW8nbVdhITJpECJtUzE+pDoof4oDdnKEJYXECqh7QHS96Tk4+JQE7dPuxck
ARJr1f0RTkAdVPFbO1OairCor2aL0QBSSStvdOtGjoFvoG+Xa7cB1b2UsPh2aeZs
M27JDWlSUUF56guJh3CnF4qoyTeF6/vbBZSsxLJs9XzpE77a/ET3HfYGUgLtOGZz
rgYCI0jETrUgndy8iiaivV/L9CLEZeLtDAYItsYRfKddyx9QMp5h1m1Pc4Eak7Bi
rtQ8ygDlcpiGR1dqe8nEJWJWCe/BSip+6Ky3rSQHlpgkkDLUiTcp/gMVS3IIwZ7a
n3jAU+lNftAIijRZA8rvNkGroVBWYkC6LVsgBF000U0fyPed7uivGFQa3/1fgR7P
RHQtbiFBxOq7yzU3WlHgaiACICPcAOmLOfgNHVy/4Qgh554+gyIYQDsLcZ4lRCAM
8HrgV+Yu7QZszs0oOuLz9+sNihL0svdTC4HogHWSTopzBu4UGlHnlVQr8tlaHb8/
wlqR56ZQG3xad/Pp8NVwmi1gUFmmfkREKzJuhMkKdT8vAO5e94hMCmIxGuFW/yR5
kEG1+7LJ5bA6opLT03hu7Vasf+EPP9eX5aUsKM9BQE8ZAEpMHQjhngW20xYgcAn/
9Q5Frfjaqi7wVT+LIh6nKDxbpMjydJatPrePGrEkUxMdV2j+Sl/DJU3Sg7OfA5k0
UYlsHnYO36Mkec4b3qN0770XgVh6TyO8QTZLlmu59vuwW3f0byi1boIFH2FwkvIl
0/ZU5tRysrU9FiJe8tLnn/isr0vd86iMXVrJlraGU9183JIWLwx8vRm7WSqNS/Qk
E2i4HscOefGrgEKSvqnLN9HzRNHP9Nqd2YEdclLoqDobMOOCDfoyGiIlrBnK2qn/
TXqAyzlhOwrdeUWPrPWPxId9Qo2YWkVfmag76o6iKQI68qMyTVhVkjM9JmzP3DrL
3m+FspGx2blKB7sx22mwgQtbGWR2Rm/f0IEhh7nIzC52XaKQCzssI1ZdrBudY4Fk
xPu3+Dlvg3Vm4E4Te8HjnOANpVjelRhC+BgO7ly26MMCFldqynkd48lo82NFHH1P
BHhm+c/H7bn8E7l24eVlSluoezD76IX0ZJrObCltz5HMHLQOgSwllV17XMZz3MTW
qm7PREYkqYJZ5V2k5Tb5UKc8Ib/X7sAbUwmCyDLy2KSqNuP8EcvU8eJ+C5MIXjZW
Z5z6OOo7FIMtV+Dzqr6oyNYRqK33V4UZTvtdeqgM98/z29M0h2rAdV7kmGXOLXwy
8R+Wns++LfBIqez2WCZqehW9Fq9AdGwMhQzlKFb4etuhH580E6PTXz/J+v8NNxlk
9ZWe/SQ42cobO0I9brrfhn92ZfsuH16fFA8MMHP/9x3P7XF3V/AKehPk4ppPbduK
bZ20PronZvNei2J0fkSyi4nIawUHLOZZB3CK3qJY1CIFXku4sEUJzKv6fZwwnVUR
Oq9yKYJIg61fYeHL8p/mjgzIPTsQDAlETu7/RSDVBZzeFlPv+e1MwfBeCAzEF6LW
zd3ZYkN3H0FMcPaesC5ZWZagSxz7S7JYJTNjsEgkuzhY0hRY6dD2K9M1izWz4uhK
eQuA+AvPUlaqcooAjNq5qCHhRtJ1SrLP0NlpVmyabpoxahgoE3597848l+VTX3sx
j0Ai+dUpIC92Evv/S+xhQ8tkRWvagXlFdcloaBhh121aVxERXpm4KmOpG7c7nd+O
sMQSB0HvRJebBggWnzDNBqzjwlY62jQxbaSs2mihVK6lHTvxYh26xN8SQ2gcjKOw
1J8MF9pyFcaDn3Mf5ryNkNcJGAIJB0LzT1IrB2s0tc/Rv6o6tL4HWYosCNzTv9iA
a+eyx++k4mboFZWAk4Z4pWosAKsd3xf2we+ZFwl4RRQ06e3dkJrsbkTZQhGR8vT+
NCk/S0nWQ2LkgMXGAHU3TLY8BG3qR5GpBYnEjUPeIU9J0WZJUvkLPQRdhWUtk11o
iHClLveTuBZqt4ZIjo8GH6jhKw2kZErSufU487Ugkoam4HNT7XoT5rVsBje3cX37
dxH5HtUf9fbhHY46ggJhPjcT5X7WocHK39oY1s4uxfPZDWJIXPiTKjEQlsewq4ee
XcahwpEhMI/87pDjyYChy7awMP1V4YyTo1kJAyyDWBz1LgadEqWQdRmlfnVpdeJX
8wAWOzstdTfNpB7Eo7zq8KeC3xsr3TGeOFEkA0IlcMfgf6PGVu7ZMeNGpcGpW+eu
BCEEN8UOGj+oiaukwJMx1ExpwOGLB7l1UR1Znu2Q0qgKJXghthK8X8Z4zwzK3XRI
/YnwA4voPNSe/nQMgzfEC4jObLxkT53zFTDdghMUcaOdiqfy3LTo7Xf4Hf2CovHh
v2ZRgajf2R9G2j0OLJ9+iRiwHy6AzKFryTDCTvCz3h2zsVyL4KXV6zDVyewjsV0a
63THqI7W4DMT/cmaEj+eYVR6YgRY2iXFeVjaVtyWFuvqOmKA5lSul6Qktu8Lr5DX
3yys04tR08e0ba9F1QKTQBDIGZ058DmewWZZhZV7HLlXC94IrFnhQsnfT4IBh/Ve
oojSHF6MTl6HaLlwY9hJ9dHR4/tps/vVB3Dh/p9TclpBqxwBB1ijCJzhdFR2WUss
VxxN8fL7PMRCz1ya7MGcgvjPmawZL7p2J2LJNxy9aC0IDJl4u/0imRio8PJ+xpEo
VELwDnOlN2pLmWBiIIcKQUQZsETVrTp0NaYDqb9fkz+w7HN66eMpWy94f2HaiRtB
1HJMMWQq1B1aObxK3ardL86lKHWSWxuFNIevuZ+EvWZ+c3Oov4IGbQE4vLcTg8++
D15osRfRjMAa8IlsCZC7N7Nvfs/0n4YT6Ar1IbQCV8qTqlmIT+3MnnHz8e9mGnPW
y9mu8mjrsCFwWWudF4czLoNVgTKBnVdQWtTEXGNZ2XI04wmtYZZBqp3+rrAyavMO
2gHBdcEWrhYyTIcNxfr4MfjM47MrYTB9iMEmLHPEuoYRZSd7qbRyckiRZuJqep8m
jkp+gGtnjeeYm5dkW1Ddorazqta0nXrAFaUDVmiApUOSJH3Le0aZRp7mj/o94RoH
F6ettSNjzMgfUYMSLVYOef8IxvNEEOFy96ktwR3cBrT9ptR+IyDromFNxi550f9T
BR8JJFSJTdGRHTat6afFKaVhbmW7muOMLeENwUEQZmjhL9i3x8bZieHAXa7cXTxY
hfXgaSjenoYfePV2TLPU56Jxzl0JtGx4Z6HSsBMo9vk6dSdzIN8dI8OVPlI/DA4w
uEp8Fz0KdwFxFg3AP6Fc0vZpO5XlDgLZCeCvmeE/koSCgW1kkqvGMd/rogtTftQl
FeiLsRS9Yw3mpbzVYMKpO8iEr874/NSgWXLVkNaTtOXimcDrpKQzNKjr4dtt3ELn
QjiigAfWSIVBF9UE7TxJCnssWT7fhUJUNX2AiQwbPGZ+2tggxKQREAN1Ez5/5Ruv
mZ5EOgKz8acZkp0+WbhaqdCnwrNiFigy7EtpXwT31G0zzgLbZrlvPqOmrOs/4iYA
R3T1wSy3AM9oYIcJ7z9pUEQGuUs9vfAh7cySf0T+UjC4tgkIsDHVPSP26+2BBmB5
2VR8luai859xlK86p+MtPvBVkQQgribG6A6XnIT9BsEKZmVGwokYmQOMyR7sEcig
wt1/Hr49m9fMboxehK4oq17+nRklOsj/CHLICjB9qHJYoLnqD/zMV24axKvp0ra/
hTmEvxHEn1L+yc6GZxXA+6EVlEFvQyOiG7IFwmb815SOXpJgh+Bk2YdxIzZVHxKA
ReVUyGlBHLVSSiFBpOOw0LzxAu5QHuTRIKJRdFUOzLOyQLE5x4GMgZfJ0EnJWeDF
ExuR4t2+IyyoSR6Yy7hCqapDruYzNiV/Jem6iMidTDfLJPwhcu7hkut1spOz9/LV
KQfVbSEna1ScG/IaZ5dtFw1+jgIQ5EeZ4pyves6M5oM3yTsPyvI55cxIMY1zLBSY
duqb3B9VaQnfCAU1TuQF6ZpBIQ5rgmmEuqY5l18sEi0Oz4rhR2+PaqhyL4MHJBGz
B55Npehr+HGLSGLWl3jj5t5g00cH/1siLelxaZsloS+/4sC7wdvgFX2qKIcUv9nc
cO6Kcl66lDXgtPit+8kQJEd6YwfMKYfH0hM9JhGp+xSIAj1BP/InQyoVE+dlhgr4
slzHv+2fD0lvBmOp0xzyFvtQivjucqTJNhqU4ZBLfrkySLb3jp5D95+afGMn7xma
TbYsXzNf61Cjq3c7JKtkS3nXAg3FN1LedZHKqETLF6rMhCZD1CnLzl/4+waXxfx3
t9Y7XsIRH7TjpRiL0v8worFk6iACF3jxyNuFdXEIlKMZ+Hl1Esui1pqYD6tgT2cF
BrHmjXqGlL4SeeDWjULKg6hmEt9iNtAicE06Pay3M73bcFX2h7fkL3BlKASnAd1k

//pragma protect end_data_block
//pragma protect digest_block
zhgy0EMXDNkO58WETA3QUPkpd4w=
//pragma protect end_digest_block
//pragma protect end_protected
